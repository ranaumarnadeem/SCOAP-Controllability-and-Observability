module s15850(CK, g100, g101, g102, g103, g10377, g10379, g104, g10455,
     g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109,
     g11163, g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185,
     g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700, g1712,
     g18, g1957, g1960, g1961, g23, g2355, g2601, g2602, g2603, g2604,
     g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648,
     g27, g28, g29, g2986, g30, g3007, g3069, g31, g3327, g41, g4171,
     g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180,
     g4181, g4191, g4192, g4193, g4194, g4195, g4196, g4197, g4198,
     g4199, g42, g4200, g4201, g4202, g4203, g4204, g4205, g4206,
     g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214, g4215,
     g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, g5105,
     g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258,
     g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267,
     g6268, g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276,
     g6277, g6278, g6279, g6280, g6281, g6282, g6283, g6284, g6285,
     g6842, g6920, g6926, g6932, g6942, g6949, g6955, g741, g742, g743,
     g744, g750, g7744, g8061, g8062, g82, g8271, g83, g8313, g8316,
     g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352,
     g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
     g872, g873, g877, g88, g881, g886, g889, g89, g892, g895, g8976,
     g8977, g8978, g8979, g898, g8980, g8981, g8982, g8983, g8984,
     g8985, g8986, g90, g901, g904, g907, g91, g910, g913, g916, g919,
     g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, SE,
     scan_in, scan_out, dft_sdi_1, dft_sdo_1, dft_sdi_2, dft_sdo_2,
     dft_sdi_3, dft_sdo_3, dft_sdi_4, dft_sdo_4, dft_sdi_5, dft_sdo_5,
     dft_sdi_6, dft_sdo_6, dft_sdi_7, dft_sdo_7, dft_sdi_8, dft_sdo_8,
     dft_sdi_9, dft_sdo_9, dft_sdi_10, dft_sdo_10, dft_sdi_11,
     dft_sdo_11, dft_sdi_12, dft_sdo_12, dft_sdi_13, dft_sdo_13,
     dft_sdi_14, dft_sdo_14, dft_sdi_15, dft_sdo_15, dft_sdi_16,
     dft_sdo_16, dft_sdi_17, dft_sdo_17, dft_sdi_18, dft_sdo_18,
     dft_sdi_19, dft_sdo_19, dft_sdi_20, dft_sdo_20, dft_sdi_21,
     dft_sdo_21, dft_sdi_22, dft_sdo_22, dft_sdi_23, dft_sdo_23,
     dft_sdi_24, dft_sdo_24, dft_sdi_25, dft_sdo_25, dft_sdi_26,
     dft_sdo_26, dft_sdi_27, dft_sdo_27, dft_sdi_28, dft_sdo_28,
     dft_sdi_29, dft_sdo_29);
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176,
       g1179, g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203,
       g1696, g1700, g1712, g18, g1960, g1961, g23, g27, g28, g29, g30,
       g31, g41, g42, g43, g44, g45, g46, g47, g48, g741, g742, g743,
       g744, g750, g82, g83, g84, g85, g86, g87, g872, g873, g877, g88,
       g881, g886, g889, g89, g892, g895, g898, g90, g901, g904, g907,
       g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g95,
       g96, g99, SE, scan_in, dft_sdi_1, dft_sdi_2, dft_sdi_3,
       dft_sdi_4, dft_sdi_5, dft_sdi_6, dft_sdi_7, dft_sdi_8,
       dft_sdi_9, dft_sdi_10, dft_sdi_11, dft_sdi_12, dft_sdi_13,
       dft_sdi_14, dft_sdi_15, dft_sdi_16, dft_sdi_17, dft_sdi_18,
       dft_sdi_19, dft_sdi_20, dft_sdi_21, dft_sdi_22, dft_sdi_23,
       dft_sdi_24, dft_sdi_25, dft_sdi_26, dft_sdi_27, dft_sdi_28,
       dft_sdi_29;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463,
       g10465, g10628, g10801, g11163, g11206, g11489, g1957, g2355,
       g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609,
       g2610, g2611, g2612, g2648, g2986, g3007, g3069, g3327, g4171,
       g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180,
       g4181, g4191, g4192, g4193, g4194, g4195, g4196, g4197, g4198,
       g4199, g4200, g4201, g4202, g4203, g4204, g4205, g4206, g4207,
       g4208, g4209, g4210, g4211, g4212, g4213, g4214, g4215, g4216,
       g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253, g6254,
       g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
       g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272,
       g6273, g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281,
       g6282, g6283, g6284, g6285, g6842, g6920, g6926, g6932, g6942,
       g6949, g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318,
       g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561,
       g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979,
       g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961,
       scan_out, dft_sdo_1, dft_sdo_2, dft_sdo_3, dft_sdo_4, dft_sdo_5,
       dft_sdo_6, dft_sdo_7, dft_sdo_8, dft_sdo_9, dft_sdo_10,
       dft_sdo_11, dft_sdo_12, dft_sdo_13, dft_sdo_14, dft_sdo_15,
       dft_sdo_16, dft_sdo_17, dft_sdo_18, dft_sdo_19, dft_sdo_20,
       dft_sdo_21, dft_sdo_22, dft_sdo_23, dft_sdo_24, dft_sdo_25,
       dft_sdo_26, dft_sdo_27, dft_sdo_28, dft_sdo_29;
  wire CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176,
       g1179, g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203,
       g1696, g1700, g1712, g18, g1960, g1961, g23, g27, g28, g29, g30,
       g31, g41, g42, g43, g44, g45, g46, g47, g48, g741, g742, g743,
       g744, g750, g82, g83, g84, g85, g86, g87, g872, g873, g877, g88,
       g881, g886, g889, g89, g892, g895, g898, g90, g901, g904, g907,
       g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g95,
       g96, g99, SE, scan_in, dft_sdi_1, dft_sdi_2, dft_sdi_3,
       dft_sdi_4, dft_sdi_5, dft_sdi_6, dft_sdi_7, dft_sdi_8,
       dft_sdi_9, dft_sdi_10, dft_sdi_11, dft_sdi_12, dft_sdi_13,
       dft_sdi_14, dft_sdi_15, dft_sdi_16, dft_sdi_17, dft_sdi_18,
       dft_sdi_19, dft_sdi_20, dft_sdi_21, dft_sdi_22, dft_sdi_23,
       dft_sdi_24, dft_sdi_25, dft_sdi_26, dft_sdi_27, dft_sdi_28,
       dft_sdi_29;
  wire g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
       g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601,
       g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610,
       g2611, g2612, g2648, g2986, g3007, g3069, g3327, g4171, g4172,
       g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181,
       g4191, g4192, g4193, g4194, g4195, g4196, g4197, g4198, g4199,
       g4200, g4201, g4202, g4203, g4204, g4205, g4206, g4207, g4208,
       g4209, g4210, g4211, g4212, g4213, g4214, g4215, g4216, g4887,
       g4888, g5101, g5105, g5658, g5659, g5816, g6253, g6254, g6255,
       g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263, g6264,
       g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
       g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282,
       g6283, g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949,
       g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323,
       g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561, g8562,
       g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979, g8980,
       g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961,
       scan_out, dft_sdo_1, dft_sdo_2, dft_sdo_3, dft_sdo_4, dft_sdo_5,
       dft_sdo_6, dft_sdo_7, dft_sdo_8, dft_sdo_9, dft_sdo_10,
       dft_sdo_11, dft_sdo_12, dft_sdo_13, dft_sdo_14, dft_sdo_15,
       dft_sdo_16, dft_sdo_17, dft_sdo_18, dft_sdo_19, dft_sdo_20,
       dft_sdo_21, dft_sdo_22, dft_sdo_23, dft_sdo_24, dft_sdo_25,
       dft_sdo_26, dft_sdo_27, dft_sdo_28, dft_sdo_29;
  wire UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2,
       UNCONNECTED3, UNCONNECTED4, UNCONNECTED5, UNCONNECTED6;
  wire UNCONNECTED7, UNCONNECTED8, UNCONNECTED9, UNCONNECTED10,
       UNCONNECTED11, UNCONNECTED12, UNCONNECTED13, UNCONNECTED14;
  wire UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18,
       UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22;
  wire UNCONNECTED23, UNCONNECTED24, UNCONNECTED25, UNCONNECTED26,
       UNCONNECTED27, UNCONNECTED28, UNCONNECTED29, UNCONNECTED30;
  wire UNCONNECTED31, UNCONNECTED32, UNCONNECTED33, UNCONNECTED34,
       UNCONNECTED35, UNCONNECTED36, UNCONNECTED37, UNCONNECTED38;
  wire UNCONNECTED39, UNCONNECTED40, UNCONNECTED41, UNCONNECTED42,
       UNCONNECTED43, UNCONNECTED44, UNCONNECTED45, UNCONNECTED46;
  wire UNCONNECTED47, g1, g4, g7, g8, g9, g16, g17;
  wire g32, g33, g34, g35, g36, g37, g38, g39;
  wire g40, g105, g108, g115, g123, g127, g131, g135;
  wire g139, g143, g148, g153, g158, g162, g166, g170;
  wire g174, g178, g182, g186, g192, g197, g201, g207;
  wire g213, g219, g225, g231, g237, g243, g248, g253;
  wire g254, g255, g256, g257, g258, g259, g260, g261;
  wire g262, g263, g266, g269, g272, g275, g278, g281;
  wire g284, g287, g290, g293, g296, g299, g302, g305;
  wire g309, g312, g315, g318, g321, g324, g327, g330;
  wire g333, g336, g339, g342, g345, g348, g351, g354;
  wire g357, g360, g363, g366, g369, g374, g378, g382;
  wire g386, g391, g396, g401, g406, g411, g416, g421;
  wire g426, g431, g435, g440, g444, g448, g452, g456;
  wire g461, g466, g471, g476, g481, g486, g491, g496;
  wire g501, g506, g511, g516, g521, g525, g530, g534;
  wire g538, g542, g546, g549, g554, g557, g560, g563;
  wire g566, g569, g572, g575, g590, g591, g599, g605;
  wire g611, g617, g622, g627, g630, g631, g632, g635;
  wire g636, g639, g643, g646, g650, g654, g658, g664;
  wire g668, g673, g677, g682, g686, g691, g695, g700;
  wire g704, g709, g713, g718, g722, g727, g731, g736;
  wire g745, g755, g756, g757, g794, g798, g802, g806;
  wire g810, g814, g818, g822, g826, g829, g833, g837;
  wire g841, g845, g849, g853, g857, g861, g868, g869;
  wire g874, g875, g876, g944, g947, g950, g953, g956;
  wire g959, g962, g965, g968, g971, g976, g981, g986;
  wire g991, g995, g999, g1003, g1007, g1011, g1015, g1019;
  wire g1023, g1027, g1032, g1068, g1071, g1074, g1077, g1080;
  wire g1083, g1086, g1089, g1092, g1095, g1098, g1212, g1217;
  wire g1218, g1223, g1227, g1231, g1235, g1240, g1245, g1250;
  wire g1255, g1260, g1265, g1270, g1280, g1284, g1292, g1296;
  wire g1300, g1304, g1308, g1311, g1314, g1317, g1318, g1321;
  wire g1324, g1327, g1330, g1333, g1336, g1341, g1346, g1351;
  wire g1356, g1361, g1362, g1365, g1368, g1371, g1374, g1377;
  wire g1380, g1383, g1386, g1389, g1393, g1394, g1397, g1400;
  wire g1403, g1407, g1411, g1415, g1419, g1424, g1428, g1432;
  wire g1436, g1440, g1444, g1448, g1453, g1462, g1466, g1470;
  wire g1474, g1478, g1482, g1486, g1490, g1494, g1499, g1504;
  wire g1508, g1515, g1520, g1524, g1528, g1531, g1534, g1537;
  wire g1540, g1543, g1546, g1549, g1552, g1555, g1558, g1561;
  wire g1564, g1567, g1571, g1574, g1577, g1580, g1583, g1586;
  wire g1589, g1592, g1595, g1598, g1601, g1604, g1607, g1615;
  wire g1618, g1621, g1624, g1627, g1630, g1633, g1636, g1654;
  wire g1657, g1660, g1663, g1666, g1690, g1703, g1707, g1710;
  wire g1713, g1718, g1721, g1724, g1727, g1730, g1733, g1766;
  wire g1771, g1776, g1781, g1786, g1791, g1796, g1801, g1806;
  wire g1811, g1814, g1822, g1828, g1834, g1840, g1845, g1848;
  wire g1849, g1850, g1853, g1854, g1857, g1861, g1864, g1868;
  wire g1872, g1878, g1882, g1887, g1891, g1896, g1900, g1905;
  wire g1909, g1914, g1918, g1923, g1927, g1932, g1936, g1941;
  wire g1945, g1950, g1958, g1959, n_0, n_1, n_2, n_3;
  wire n_4, n_5, n_7, n_8, n_9, n_10, n_11, n_12;
  wire n_13, n_14, n_15, n_16, n_17, n_18, n_20, n_21;
  wire n_22, n_23, n_25, n_26, n_27, n_28, n_29, n_30;
  wire n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38;
  wire n_39, n_40, n_42, n_44, n_45, n_46, n_47, n_48;
  wire n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_67, n_68, n_69, n_70, n_71, n_72, n_73;
  wire n_74, n_75, n_76, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_88, n_89, n_90;
  wire n_91, n_92, n_94, n_95, n_96, n_97, n_98, n_99;
  wire n_100, n_101, n_102, n_103, n_104, n_105, n_106, n_107;
  wire n_108, n_109, n_111, n_112, n_113, n_115, n_116, n_117;
  wire n_118, n_119, n_121, n_122, n_123, n_124, n_125, n_126;
  wire n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134;
  wire n_135, n_136, n_137, n_139, n_140, n_142, n_143, n_144;
  wire n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152;
  wire n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160;
  wire n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168;
  wire n_169, n_170, n_171, n_172, n_174, n_175, n_176, n_177;
  wire n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185;
  wire n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193;
  wire n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_202;
  wire n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210;
  wire n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218;
  wire n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226;
  wire n_227, n_228, n_229, n_230, n_231, n_232, n_234, n_235;
  wire n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243;
  wire n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251;
  wire n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_259;
  wire n_260, n_261, n_262, n_263, n_264, n_265, n_266, n_267;
  wire n_268, n_269, n_270, n_271, n_272, n_274, n_275, n_276;
  wire n_278, n_279, n_280, n_281, n_282, n_283, n_284, n_286;
  wire n_288, n_289, n_290, n_291, n_292, n_293, n_294, n_295;
  wire n_296, n_297, n_298, n_299, n_300, n_301, n_302, n_303;
  wire n_304, n_305, n_308, n_310, n_311, n_312, n_313, n_314;
  wire n_315, n_316, n_317, n_318, n_319, n_320, n_321, n_322;
  wire n_323, n_325, n_326, n_327, n_329, n_330, n_331, n_332;
  wire n_333, n_334, n_336, n_337, n_338, n_339, n_340, n_341;
  wire n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_350;
  wire n_351, n_352, n_353, n_354, n_355, n_356, n_357, n_358;
  wire n_359, n_360, n_361, n_362, n_363, n_364, n_365, n_366;
  wire n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374;
  wire n_375, n_377, n_378, n_379, n_380, n_381, n_382, n_383;
  wire n_384, n_385, n_386, n_387, n_388, n_389, n_390, n_391;
  wire n_392, n_393, n_394, n_395, n_396, n_397, n_398, n_399;
  wire n_400, n_401, n_402, n_404, n_405, n_406, n_407, n_408;
  wire n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416;
  wire n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424;
  wire n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432;
  wire n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440;
  wire n_441, n_442, n_443, n_444, n_446, n_447, n_448, n_449;
  wire n_450, n_451, n_452, n_453, n_455, n_456, n_457, n_458;
  wire n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466;
  wire n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474;
  wire n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482;
  wire n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490;
  wire n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498;
  wire n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506;
  wire n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514;
  wire n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522;
  wire n_523, n_524, n_525, n_526, n_527, n_528, n_529, n_530;
  wire n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538;
  wire n_539, n_540, n_541, n_542, n_543, n_544, n_545, n_546;
  wire n_547, n_548, n_549, n_550, n_551, n_552, n_553, n_554;
  wire n_555, n_556, n_557, n_558, n_559, n_560, n_561, n_562;
  wire n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570;
  wire n_571, n_572, n_573, n_574, n_575, n_576, n_577, n_578;
  wire n_579, n_580, n_581, n_582, n_583, n_584, n_585, n_586;
  wire n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594;
  wire n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602;
  wire n_603, n_604, n_605, n_606, n_607, n_608, n_609, n_610;
  wire n_611, n_612, n_613, n_614, n_615, n_616, n_617, n_618;
  wire n_619, n_620, n_621, n_622, n_623, n_624, n_625, n_626;
  wire n_627, n_628, n_629, n_630, n_631, n_632, n_633, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659;
  wire n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667;
  wire n_668, n_669, n_670, n_671, n_672, n_673, n_674, n_675;
  wire n_676, n_677, n_678, n_679, n_680, n_681, n_682, n_683;
  wire n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691;
  wire n_692, n_693, n_694, n_695, n_696, n_697, n_698, n_699;
  wire n_700, n_701, n_702, n_703, n_704, n_705, n_706, n_707;
  wire n_708, n_709, n_710, n_711, n_712, n_713, n_714, n_715;
  wire n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723;
  wire n_724, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_737, n_738, n_739;
  wire n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747;
  wire n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755;
  wire n_756, n_757, n_758, n_759, n_760, n_761, n_762, n_763;
  wire n_764, n_765, n_766, n_767, n_768, n_769, n_770, n_771;
  wire n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779;
  wire n_780, n_781, n_782, n_783, n_784, n_785, n_786, n_787;
  wire n_788, n_789, n_790, n_791, n_792, n_793, n_794, n_795;
  wire n_796, n_797, n_798, n_799, n_800, n_801, n_802, n_803;
  wire n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811;
  wire n_812, n_813, n_814, n_815, n_816, n_817, n_818, n_819;
  wire n_820, n_821, n_822, n_823, n_824, n_825, n_826, n_827;
  wire n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835;
  wire n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843;
  wire n_844, n_845, n_846, n_847, n_848, n_849, n_850, n_851;
  wire n_852, n_853, n_854, n_855, n_856, n_857, n_858, n_859;
  wire n_860, n_861, n_862, n_864, n_865, n_866, n_867, n_868;
  wire n_869, n_870, n_871, n_873, n_874, n_875, n_876, n_877;
  wire n_878, n_879, n_880, n_881, n_882, n_883, n_884, n_885;
  wire n_886, n_887, n_888, n_889, n_890, n_891, n_892, n_893;
  wire n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901;
  wire n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909;
  wire n_910, n_911, n_912, n_913, n_914, n_915, n_916, n_917;
  wire n_918, n_919, n_920, n_921, n_922, n_923, n_924, n_925;
  wire n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933;
  wire n_934, n_935, n_936, n_937, n_938, n_939, n_940, n_941;
  wire n_942, n_943, n_944, n_945, n_946, n_947, n_948, n_949;
  wire n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957;
  wire n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965;
  wire n_966, n_967, n_968, n_969, n_970, n_971, n_972, n_973;
  wire n_974, n_975, n_976, n_977, n_978, n_979, n_980, n_981;
  wire n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989;
  wire n_990, n_991, n_992, n_993, n_994, n_995, n_996, n_997;
  wire n_998, n_999, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005;
  wire n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013;
  wire n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021;
  wire n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029;
  wire n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037;
  wire n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045;
  wire n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053;
  wire n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061;
  wire n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069;
  wire n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077;
  wire n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085;
  wire n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093;
  wire n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101;
  wire n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109;
  wire n_1110, n_1111, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118;
  wire n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126;
  wire n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134;
  wire n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142;
  wire n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150;
  wire n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158;
  wire n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1167;
  wire n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175;
  wire n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183;
  wire n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223;
  wire n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231;
  wire n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239;
  wire n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247;
  wire n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256;
  wire n_1257, n_1258, n_1259, n_1260, n_1263, n_1264, n_1265, n_1266;
  wire n_1267, n_1268, n_1270, n_1271, n_1273, n_1274, n_1275, n_1276;
  wire n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284;
  wire n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292;
  wire n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300;
  wire n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1308, n_1309;
  wire n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317;
  wire n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1325, n_1327;
  wire n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335;
  wire n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343;
  wire n_1344, n_1345, n_1346, n_1347, n_1348, n_1350, n_1351, n_1353;
  wire n_1354, n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361;
  wire n_1362, n_1363, n_1364, n_1365, n_1366, n_1368, n_1369, n_1370;
  wire n_1372, n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379;
  wire n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, n_1387, n_1388;
  wire n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, n_1396, n_1397;
  wire n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405;
  wire n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413;
  wire n_1414, n_1415, n_1416, n_1418, n_1419, n_1420, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430;
  wire n_1431, n_1432, n_1433, n_1435, n_1436, n_1437, n_1438, n_1439;
  wire n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1447, n_1448;
  wire n_1449, n_1451, n_1452, n_1453, n_1454, n_1455, n_1457, n_1458;
  wire n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466;
  wire n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1484;
  wire n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492;
  wire n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500;
  wire n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508;
  wire n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516;
  wire n_1517, n_1518, n_1519, n_1520, n_1522, n_1523, n_1524, n_1525;
  wire n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533;
  wire n_1534, n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541;
  wire n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549;
  wire n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, n_1557;
  wire n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565;
  wire n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573;
  wire n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582;
  wire n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1590, n_1591;
  wire n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
  wire n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607;
  wire n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615;
  wire n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623;
  wire n_1624, n_1625, n_1626, n_1627, n_1628, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1640, n_1641;
  wire n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649;
  wire n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1657, n_1658;
  wire n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667;
  wire n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676;
  wire n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684;
  wire n_1685, n_1686, n_1687, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702;
  wire n_1703, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712;
  wire n_1713, n_1714, n_1715, n_1731, n_1732, n_1733, n_1734, n_1735;
  wire n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742;
  assign g9961 = g9451;
  assign g8986 = 1'b0;
  assign g8985 = 1'b0;
  assign g8984 = 1'b1;
  assign g8983 = 1'b0;
  assign g8982 = 1'b1;
  assign g8981 = 1'b0;
  assign g8980 = 1'b1;
  assign g8979 = 1'b0;
  assign g8978 = 1'b1;
  assign g8977 = 1'b0;
  assign g8976 = 1'b1;
  assign g8566 = g6955;
  assign g8565 = g6949;
  assign g8564 = g6942;
  assign g8563 = g6932;
  assign g8562 = g6926;
  assign g8561 = g6920;
  assign g8352 = g82;
  assign g8349 = g82;
  assign g8347 = 1'b1;
  assign g8340 = 1'b1;
  assign g8335 = g82;
  assign g8331 = 1'b1;
  assign g8328 = g82;
  assign g8323 = 1'b1;
  assign g8318 = g82;
  assign g8316 = 1'b1;
  assign g8313 = g82;
  assign g8271 = g5816;
  assign g8062 = g873;
  assign g8061 = g872;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6284 = g104;
  assign g6283 = g103;
  assign g6282 = g102;
  assign g6281 = g101;
  assign g6280 = g100;
  assign g6279 = g99;
  assign g6278 = g96;
  assign g6277 = g95;
  assign g6276 = g94;
  assign g6275 = g93;
  assign g6274 = g92;
  assign g6273 = g91;
  assign g6272 = g90;
  assign g6271 = g89;
  assign g6270 = g88;
  assign g6269 = g87;
  assign g6268 = g86;
  assign g6267 = g85;
  assign g6266 = g84;
  assign g6265 = g83;
  assign g6264 = g82;
  assign g6263 = g48;
  assign g6262 = g47;
  assign g6261 = g46;
  assign g6260 = g45;
  assign g6259 = g44;
  assign g6258 = g43;
  assign g6257 = g42;
  assign g6256 = g41;
  assign g6255 = g31;
  assign g6254 = g30;
  assign g6253 = g29;
  assign g5105 = g873;
  assign g5101 = g872;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g4216 = g1194;
  assign g4215 = g1191;
  assign g4214 = g1188;
  assign g4213 = g1185;
  assign g4212 = g1182;
  assign g4211 = g1179;
  assign g4210 = g1176;
  assign g4209 = g1173;
  assign g4208 = g1203;
  assign g4207 = g1200;
  assign g4206 = g1197;
  assign g4205 = g1170;
  assign g4204 = g922;
  assign g4203 = g919;
  assign g4202 = g916;
  assign g4201 = g913;
  assign g4200 = g910;
  assign g4199 = g907;
  assign g4198 = g904;
  assign g4197 = g901;
  assign g4196 = g925;
  assign g4195 = g898;
  assign g4194 = g895;
  assign g4193 = g892;
  assign g4192 = g889;
  assign g4191 = g886;
  assign g2986 = 1'b0;
  assign g2612 = g2606;
  assign g2611 = g2605;
  assign g2610 = g2601;
  assign g2609 = g2604;
  assign g2608 = g2603;
  assign g2607 = g2602;
  assign g2355 = g18;
  assign g11489 = 1'b0;
  SDFFX1 DFF_317_Q_reg(.CK (CK), .D (n_1708), .SI (n_200), .SE (SE), .Q
       (g953), .QN (n_384));
  SDFFX1 DFF_312_Q_reg(.CK (CK), .D (n_1706), .SI (n_262), .SE (SE), .Q
       (g944), .QN (n_383));
  SDFFX1 DFF_454_Q_reg(.CK (CK), .D (n_1709), .SI (n_247), .SE (SE), .Q
       (g947), .QN (n_382));
  SDFFX1 DFF_365_Q_reg(.CK (CK), .D (n_1715), .SI (g182), .SE (SE), .Q
       (g950), .QN (n_381));
  SDFFX1 DFF_106_Q_reg(.CK (CK), .D (n_1712), .SI (n_352), .SE (SE), .Q
       (g959), .QN (n_380));
  SDFFX1 DFF_408_Q_reg(.CK (CK), .D (n_1711), .SI (n_63), .SE (SE), .Q
       (g956), .QN (n_379));
  SDFFX1 DFF_351_Q_reg(.CK (CK), .D (n_1714), .SI (n_228), .SE (SE), .Q
       (g968), .QN (n_378));
  SDFFX1 DFF_148_Q_reg(.CK (CK), .D (n_1710), .SI (n_353), .SE (SE), .Q
       (g962), .QN (n_377));
  SDFFX1 DFF_181_Q_reg(.CK (CK), .D (n_1707), .SI (n_154), .SE (SE), .Q
       (g965), .QN (dft_sdo_9));
  SDFFX1 DFF_52_Q_reg(.CK (CK), .D (n_1703), .SI (n_302), .SE (SE), .Q
       (g981), .QN (n_375));
  SDFFX1 DFF_14_Q_reg(.CK (CK), .D (n_1699), .SI (n_332), .SE (SE), .Q
       (g976), .QN (n_374));
  SDFFX1 DFF_293_Q_reg(.CK (CK), .D (n_1700), .SI (n_46), .SE (SE), .Q
       (g986), .QN (n_373));
  SDFFX1 DFF_294_Q_reg(.CK (CK), .D (n_1702), .SI (n_373), .SE (SE), .Q
       (g971), .QN (n_372));
  MX2X1 g37519__2398(.A (g837), .B (g950), .S0 (n_1713), .Y (n_1715));
  MX2X1 g37518__5107(.A (g861), .B (g968), .S0 (n_1713), .Y (n_1714));
  MX2X1 g37517__6260(.A (g849), .B (g959), .S0 (n_1713), .Y (n_1712));
  MX2X1 g37520__4319(.A (g845), .B (g956), .S0 (n_1713), .Y (n_1711));
  MX2X1 g37523__8428(.A (g853), .B (g962), .S0 (n_1713), .Y (n_1710));
  MX2X1 g37522__5526(.A (g833), .B (g947), .S0 (n_1713), .Y (n_1709));
  MX2X1 g37521__6783(.A (g841), .B (g953), .S0 (n_1713), .Y (n_1708));
  MX2X1 g37524__3680(.A (g857), .B (g965), .S0 (n_1713), .Y (n_1707));
  MX2X1 g37510__1617(.A (g829), .B (g944), .S0 (n_1713), .Y (n_1706));
  AND2X2 g37528__2802(.A (n_1449), .B (g10628), .Y (g11206));
  AOI21X1 g37503__1705(.A0 (n_1693), .A1 (n_1691), .B0 (n_1701), .Y
       (n_1703));
  NOR2X1 g37525__5122(.A (n_1701), .B (n_1689), .Y (n_1702));
  NOR2X1 g37527__8246(.A (n_1701), .B (n_1695), .Y (n_1700));
  NOR2X1 g37512__7098(.A (n_1701), .B (n_1731), .Y (n_1699));
  AOI221X1 g37550__6131(.A0 (g877), .A1 (n_1407), .B0 (g109), .B1
       (n_1279), .C0 (n_1696), .Y (g10628));
  OAI21X1 g37555__1881(.A0 (n_1698), .A1 (n_1683), .B0 (n_1690), .Y
       (n_1713));
  OAI21X1 g37553__5115(.A0 (g869), .A1 (n_1697), .B0 (g109), .Y
       (n_1701));
  INVX1 g37597(.A (n_1697), .Y (n_1698));
  OAI22X1 g37563__7482(.A0 (g757), .A1 (n_1424), .B0 (n_406), .B1
       (n_1404), .Y (n_1696));
  NAND2X1 g37606__4733(.A (g757), .B (n_1278), .Y (n_1697));
  CLKXOR2X1 g37572__6161(.A (g986), .B (n_1692), .Y (n_1695));
  NAND2X1 g37599__9945(.A (g981), .B (n_1692), .Y (n_1693));
  NAND3X1 g37532__2883(.A (g976), .B (n_1686), .C (n_1687), .Y
       (n_1691));
  SDFFX1 DFF_37_Q_reg(.CK (CK), .D (n_1690), .SI (n_236), .SE (SE), .Q
       (UNCONNECTED), .QN (g757));
  SDFFX1 DFF_289_Q_reg(.CK (CK), .D (n_1684), .SI (n_198), .SE (SE), .Q
       (g1394), .QN (n_371));
  XNOR2X1 g37598__2346(.A (n_1690), .B (g971), .Y (n_1689));
  OR2X1 g37641__1666(.A (n_1686), .B (n_1685), .Y (n_1692));
  AND2X1 g37640__7410(.A (n_1690), .B (g971), .Y (n_1687));
  INVX1 g37672(.A (n_1690), .Y (n_1685));
  SDFFX1 DFF_400_Q_reg(.CK (CK), .D (n_1681), .SI (n_128), .SE (SE), .Q
       (g201), .QN (n_370));
  NOR3X1 g37674__6417(.A (n_1651), .B (n_1682), .C (n_1662), .Y
       (n_1690));
  AOI211X1 g37533__5477(.A0 (g1393), .A1 (n_394), .B0 (n_1683), .C0
       (g115), .Y (n_1684));
  SDFFX1 DFF_473_Q_reg(.CK (CK), .D (n_1680), .SI (g1710), .SE (SE), .Q
       (g115), .QN (n_369));
  SDFFX1 DFF_452_Q_reg(.CK (CK), .D (n_1679), .SI (n_199), .SE (SE), .Q
       (UNCONNECTED0), .QN (g1393));
  AOI211X1 g37723__2398(.A0 (g318), .A1 (g386), .B0 (n_1564), .C0
       (n_1676), .Y (n_1682));
  OAI21X1 g37559__5107(.A0 (n_1675), .A1 (n_1677), .B0 (n_1678), .Y
       (n_1681));
  SDFFX1 DFF_263_Q_reg(.CK (CK), .D (n_1672), .SI (n_64), .SE (SE), .Q
       (g336), .QN (n_368));
  CLKAND2X2 g37600__6260(.A (g1394), .B (n_1679), .Y (n_1680));
  OAI211X1 g37603__4319(.A0 (n_1677), .A1 (n_1674), .B0 (g109), .C0
       (n_473), .Y (n_1678));
  SDFFX1 DFF_266_Q_reg(.CK (CK), .D (n_1670), .SI (n_362), .SE (SE), .Q
       (g345), .QN (n_367));
  NAND3X1 g37729__8428(.A (n_1406), .B (n_1480), .C (n_1671), .Y
       (n_1676));
  NOR4X1 g37637__5526(.A (g1389), .B (g197), .C (n_1675), .D (n_1673),
       .Y (n_1679));
  NOR2X1 g37678__6783(.A (g197), .B (n_1673), .Y (n_1674));
  MX2X1 g37485__3680(.A (g336), .B (n_1733), .S0 (n_1669), .Y (n_1672));
  AOI211X1 g37733__1617(.A0 (g324), .A1 (g396), .B0 (n_1665), .C0
       (n_1667), .Y (n_1671));
  MX2X1 g37486__2802(.A (g345), .B (n_1666), .S0 (n_1669), .Y (n_1670));
  SDFFX1 DFF_124_Q_reg(.CK (CK), .D (n_1664), .SI (n_260), .SE (SE), .Q
       (g426), .QN (n_366));
  NAND4X1 g37681__1705(.A (g248), .B (g243), .C (g192), .D (n_1660), .Y
       (n_1673));
  OAI22X1 g37746__8246(.A0 (n_1653), .A1 (n_1657), .B0 (g318), .B1
       (g386), .Y (n_1667));
  CLKXOR2X1 g37489__7098(.A (n_1655), .B (n_1658), .Y (n_1666));
  OAI222X1 g37747__6131(.A0 (g315), .A1 (n_1661), .B0 (g305), .B1
       (n_1663), .C0 (n_1626), .C1 (g426), .Y (n_1665));
  OAI22X1 g37658__1881(.A0 (n_1663), .A1 (n_1662), .B0 (n_1661), .B1
       (n_1652), .Y (n_1664));
  NOR4X1 g37707__5115(.A (g213), .B (g1400), .C (n_1654), .D (g1374),
       .Y (n_1660));
  CLKINVX1 g37757(.A (n_1663), .Y (n_1657));
  CLKXOR2X1 g37492__7482(.A (n_1539), .B (n_1650), .Y (n_1658));
  NAND4X1 g37736__4733(.A (g1397), .B (g219), .C (n_1649), .D (n_1445),
       .Y (n_1654));
  OAI22X1 g37666__6161(.A0 (n_923), .A1 (n_1662), .B0 (n_1653), .B1
       (n_1652), .Y (n_1655));
  MX2X1 g37761__9315(.A (n_885), .B (n_1653), .S0 (n_1651), .Y
       (n_1663));
  CLKXOR2X1 g37506__9945(.A (n_1560), .B (n_1648), .Y (n_1650));
  SDFFX1 DFF_337_Q_reg(.CK (CK), .D (n_1646), .SI (g630), .SE (SE), .Q
       (g148), .QN (n_365));
  SDFFX1 DFF_34_Q_reg(.CK (CK), .D (n_1647), .SI (g243), .SE (SE), .Q
       (g1499), .QN (n_364));
  NOR4X1 g37752__2883(.A (g186), .B (g207), .C (g1377), .D (n_1645), .Y
       (n_1649));
  SDFFX1 DFF_4_Q_reg(.CK (CK), .D (n_1643), .SI (n_308), .SE (SE), .Q
       (g123), .QN (n_363));
  CLKINVX2 g37771(.A (g305), .Y (n_1653));
  CLKXOR2X1 g37760__2346(.A (g197), .B (n_1644), .Y (n_1677));
  SDFFX1 DFF_265_Q_reg(.CK (CK), .D (g253), .SI (n_327), .SE (SE), .Q
       (g305), .QN (n_362));
  SDFFX1 DFF_440_Q_reg(.CK (CK), .D (n_1638), .SI (g1490), .SE (SE), .Q
       (g348), .QN (n_361));
  SDFFX1 DFF_26_Q_reg(.CK (CK), .D (n_1642), .SI (n_25), .SE (SE), .Q
       (g546), .QN (n_360));
  CLKXOR2X1 g37536__1666(.A (n_1581), .B (n_1637), .Y (n_1648));
  SDFFX1 DFF_109_Q_reg(.CK (CK), .D (n_1635), .SI (n_54), .SE (SE), .Q
       (g1407), .QN (n_359));
  NOR2X1 g37762__7410(.A (n_1683), .B (n_1641), .Y (n_1647));
  NOR2X1 g37763__6417(.A (n_1683), .B (n_1734), .Y (n_1646));
  NAND3X1 g37779__5477(.A (g1380), .B (g1383), .C (n_1634), .Y
       (n_1645));
  SDFFX1 DFF_482_Q_reg(.CK (CK), .D (n_1632), .SI (n_279), .SE (SE), .Q
       (g1615), .QN (n_358));
  CLKXOR2X1 g37783__2398(.A (g1386), .B (g1389), .Y (n_1644));
  NOR2X1 g37696__5107(.A (n_1683), .B (n_1633), .Y (n_1643));
  OAI22X1 g37780__6260(.A0 (n_1640), .A1 (n_1586), .B0 (n_1624), .B1
       (n_1631), .Y (n_1642));
  CLKXOR2X1 g37781__4319(.A (g1494), .B (n_1640), .Y (n_1641));
  SDFFX1 DFF_397_Q_reg(.CK (CK), .D (n_1628), .SI (n_356), .SE (SE), .Q
       (g253), .QN (n_357));
  MX2X1 g37562__5526(.A (g348), .B (n_1636), .S0 (n_1669), .Y (n_1638));
  CLKXOR2X1 g37577__6783(.A (n_1608), .B (n_1636), .Y (n_1637));
  NOR2X1 g37773__3680(.A (n_1683), .B (n_1630), .Y (n_1635));
  CLKINVX1 g37792(.A (g1386), .Y (n_1634));
  AOI21X1 g37705__1617(.A0 (n_1616), .A1 (n_1625), .B0 (g123), .Y
       (n_1633));
  MX2X1 g37788__2802(.A (g1615), .B (n_1627), .S0 (n_1631), .Y
       (n_1632));
  SDFFX1 DFF_396_Q_reg(.CK (CK), .D (n_1622), .SI (n_204), .SE (SE), .Q
       (g1386), .QN (n_356));
  CLKXOR2X1 g37791__1705(.A (n_1623), .B (g1428), .Y (n_1630));
  AOI21X1 g37802__5122(.A0 (n_1595), .A1 (g1618), .B0 (n_1627), .Y
       (n_1640));
  OAI22X1 g37660__8246(.A0 (n_1626), .A1 (n_1652), .B0 (n_651), .B1
       (n_1662), .Y (n_1636));
  NOR4X1 g37725__7098(.A (n_1621), .B (g143), .C (g148), .D (g153), .Y
       (n_1625));
  OAI21X1 g37803__6131(.A0 (g18), .A1 (n_1624), .B0 (n_1623), .Y
       (n_1628));
  INVX1 g37804(.A (n_1623), .Y (n_1627));
  AND2X1 g37810__1881(.A (g109), .B (g186), .Y (n_1622));
  NAND2X1 g37809__5115(.A (g186), .B (g18), .Y (n_1623));
  SDFFX1 DFF_29_Q_reg(.CK (CK), .D (n_1620), .SI (n_194), .SE (SE), .Q
       (g4), .QN (n_355));
  INVX1 g37816(.A (g315), .Y (n_1626));
  NAND4X1 g37743__7482(.A (g127), .B (g162), .C (g135), .D (n_1619), .Y
       (n_1621));
  SDFFX1 DFF_41_Q_reg(.CK (CK), .D (g256), .SI (dft_sdi_2), .SE (SE),
       .Q (g315), .QN (n_354));
  SDFFX1 DFF_147_Q_reg(.CK (CK), .D (n_1618), .SI (dft_sdi_8), .SE
       (SE), .Q (g153), .QN (n_353));
  SDFFX1 DFF_105_Q_reg(.CK (CK), .D (n_1615), .SI (n_137), .SE (SE), .Q
       (g186), .QN (n_352));
  SDFFX1 DFF_519_Q_reg(.CK (CK), .D (n_1613), .SI (n_127), .SE (SE), .Q
       (g1494), .QN (n_351));
  SDFFX1 DFF_69_Q_reg(.CK (CK), .D (n_1611), .SI (n_31), .SE (SE), .Q
       (g554), .QN (n_350));
  SDFFX1 DFF_128_Q_reg(.CK (CK), .D (n_1612), .SI (n_181), .SE (SE), .Q
       (g1428), .QN (dft_sdo_6));
  OAI21X1 g37739__4733(.A0 (n_1683), .A1 (n_1291), .B0 (n_1617), .Y
       (n_1620));
  NOR4X1 g37768__6161(.A (g131), .B (g139), .C (g182), .D (n_1614), .Y
       (n_1619));
  SDFFX1 DFF_79_Q_reg(.CK (CK), .D (n_1609), .SI (n_29), .SE (SE), .Q
       (g351), .QN (n_348));
  SDFFX1 DFF_516_Q_reg(.CK (CK), .D (n_1607), .SI (n_47), .SE (SE), .Q
       (g1621), .QN (n_347));
  NOR2X1 g37812__9315(.A (n_1683), .B (n_1610), .Y (n_1618));
  SDFFX1 DFF_500_Q_reg(.CK (CK), .D (n_1598), .SI (n_321), .SE (SE), .Q
       (g256), .QN (n_346));
  SDFFX1 DFF_426_Q_reg(.CK (CK), .D (n_1604), .SI (n_84), .SE (SE), .Q
       (g1537), .QN (n_345));
  SDFFX1 DFF_390_Q_reg(.CK (CK), .D (n_1603), .SI (dft_sdi_22), .SE
       (SE), .Q (g275), .QN (n_344));
  NAND3X1 g37744__9945(.A (g1494), .B (n_1616), .C (n_1605), .Y
       (n_1617));
  NOR2X1 g37834__2883(.A (g1383), .B (n_1683), .Y (n_1615));
  NAND4X1 g37793__2346(.A (g178), .B (g170), .C (g166), .D (n_1596), .Y
       (n_1614));
  NOR2X1 g37811__1666(.A (n_1683), .B (n_1601), .Y (n_1613));
  NOR2X1 g37819__7410(.A (n_1683), .B (n_1600), .Y (n_1612));
  OAI211X1 g37827__6417(.A0 (n_409), .A1 (n_1631), .B0 (n_1606), .C0
       (n_1259), .Y (n_1611));
  CLKXOR2X1 g37831__5477(.A (n_1597), .B (g158), .Y (n_1610));
  MX2X1 g37561__2398(.A (g351), .B (n_1608), .S0 (n_1669), .Y (n_1609));
  OAI21X1 g37843__5107(.A0 (n_397), .A1 (n_1631), .B0 (n_1606), .Y
       (n_1607));
  SDFFX1 DFF_189_Q_reg(.CK (CK), .D (n_1594), .SI (g869), .SE (SE), .Q
       (UNCONNECTED1), .QN (g1383));
  NOR4X1 g37754__6260(.A (g1462), .B (g1490), .C (g1499), .D (n_1593),
       .Y (n_1605));
  OAI21X1 g37826__4319(.A0 (g1490), .A1 (n_1602), .B0 (n_655), .Y
       (n_1604));
  MX2X1 g37829__8428(.A (g158), .B (g275), .S0 (n_1602), .Y (n_1603));
  CLKXOR2X1 g37832__5526(.A (g1490), .B (n_1599), .Y (n_1601));
  XNOR2X1 g37846__6783(.A (n_1599), .B (g1403), .Y (n_1600));
  INVX1 g37853(.A (n_1597), .Y (n_1598));
  NOR2X1 g37844__3680(.A (g158), .B (g174), .Y (n_1596));
  NAND2X1 g37850__1617(.A (n_1599), .B (n_1631), .Y (n_1606));
  AOI21X1 g37857__2802(.A0 (n_1595), .A1 (g554), .B0 (n_1599), .Y
       (n_1597));
  OAI22X1 g37661__1705(.A0 (g318), .A1 (n_1652), .B0 (n_621), .B1
       (n_1662), .Y (n_1608));
  SDFFX1 DFF_437_Q_reg(.CK (CK), .D (n_1592), .SI (n_178), .SE (SE), .Q
       (UNCONNECTED2), .QN (g1490));
  SDFFX1 DFF_190_Q_reg(.CK (CK), .D (n_1591), .SI (g1383), .SE (SE), .Q
       (g158), .QN (n_343));
  AND2X1 g37869__5122(.A (g109), .B (g207), .Y (n_1594));
  AND2X1 g37873__8246(.A (g18), .B (g207), .Y (n_1599));
  SDFFX1 DFF_5_Q_reg(.CK (CK), .D (n_1585), .SI (n_363), .SE (SE), .Q
       (g207), .QN (n_342));
  SDFFX1 DFF_101_Q_reg(.CK (CK), .D (n_1588), .SI (n_16), .SE (SE), .Q
       (g557), .QN (n_341));
  SDFFX1 DFF_225_Q_reg(.CK (CK), .D (g257), .SI (n_153), .SE (SE), .Q
       (UNCONNECTED3), .QN (g318));
  SDFFX1 DFF_409_Q_reg(.CK (CK), .D (n_1584), .SI (n_379), .SE (SE), .Q
       (g378), .QN (n_340));
  SDFFX1 DFF_70_Q_reg(.CK (CK), .D (n_1583), .SI (n_350), .SE (SE), .Q
       (g354), .QN (n_339));
  SDFFX1 DFF_415_Q_reg(.CK (CK), .D (n_1579), .SI (n_55), .SE (SE), .Q
       (g1403), .QN (n_338));
  NAND4X1 g37790__7098(.A (g1478), .B (g1508), .C (g1482), .D (n_1582),
       .Y (n_1593));
  NOR2X1 g37868__6131(.A (n_1683), .B (n_1590), .Y (n_1592));
  NOR2X1 g37870__1881(.A (n_1683), .B (n_1735), .Y (n_1591));
  SDFFX1 DFF_374_Q_reg(.CK (CK), .D (n_1577), .SI (n_149), .SE (SE), .Q
       (g1624), .QN (n_337));
  SDFFX1 DFF_46_Q_reg(.CK (CK), .D (n_1578), .SI (n_189), .SE (SE), .Q
       (g278), .QN (n_336));
  CLKXOR2X1 g37886__5115(.A (n_1587), .B (g1486), .Y (n_1590));
  OAI22X1 g37883__4733(.A0 (n_1587), .A1 (n_1586), .B0 (n_1563), .B1
       (n_1631), .Y (n_1588));
  SDFFX1 DFF_356_Q_reg(.CK (CK), .D (n_1573), .SI (n_111), .SE (SE), .Q
       (g257), .QN (dft_sdo_19));
  NOR2X1 g37893__6161(.A (g1380), .B (n_1683), .Y (n_1585));
  SDFFX1 DFF_326_Q_reg(.CK (CK), .D (n_1572), .SI (n_278), .SE (SE), .Q
       (g1540), .QN (n_334));
  SDFFX1 DFF_207_Q_reg(.CK (CK), .D (n_1571), .SI (n_288), .SE (SE), .Q
       (g374), .QN (n_333));
  SDFFX1 DFF_12_Q_reg(.CK (CK), .D (n_1567), .SI (n_203), .SE (SE), .Q
       (g461), .QN (n_332));
  SDFFX1 DFF_255_Q_reg(.CK (CK), .D (n_1569), .SI (dft_sdi_14), .SE
       (SE), .Q (g466), .QN (n_331));
  AOI21X1 g37490__9315(.A0 (n_1529), .A1 (n_1568), .B0 (n_1570), .Y
       (n_1584));
  MX2X1 g37557__9945(.A (g354), .B (n_1580), .S0 (n_1669), .Y (n_1583));
  AND4X2 g37828__2883(.A (g1474), .B (dft_sdo_8), .C (g1466), .D
       (n_1565), .Y (n_1582));
  CLKXOR2X1 g37576__2346(.A (n_1535), .B (n_1580), .Y (n_1581));
  NOR2X1 g37875__1666(.A (n_1683), .B (n_1576), .Y (n_1579));
  SDFFX1 DFF_152_Q_reg(.CK (CK), .D (n_1561), .SI (n_293), .SE (SE), .Q
       (g471), .QN (n_330));
  OAI21X1 g37884__7410(.A0 (g162), .A1 (n_1602), .B0 (n_642), .Y
       (n_1578));
  MX2X1 g37899__6417(.A (g1624), .B (n_1575), .S0 (n_1631), .Y
       (n_1577));
  SDFFX1 DFF_487_Q_reg(.CK (CK), .D (n_1554), .SI (n_101), .SE (SE), .Q
       (UNCONNECTED4), .QN (g1380));
  SDFFX1 DFF_483_Q_reg(.CK (CK), .D (n_1559), .SI (n_358), .SE (SE), .Q
       (g382), .QN (n_329));
  CLKXOR2X1 g37900__5477(.A (n_1562), .B (g1432), .Y (n_1576));
  AOI21X1 g37903__2398(.A0 (n_1595), .A1 (g1615), .B0 (n_1575), .Y
       (n_1587));
  SDFFX1 DFF_19_Q_reg(.CK (CK), .D (n_1553), .SI (n_118), .SE (SE), .Q
       (g369), .QN (scan_out));
  SDFFX1 DFF_264_Q_reg(.CK (CK), .D (n_1550), .SI (n_368), .SE (SE), .Q
       (g456), .QN (n_327));
  MX2X1 g37881__5107(.A (g1486), .B (g1540), .S0 (n_1602), .Y (n_1572));
  NOR2X1 g37504__6260(.A (n_1570), .B (n_1555), .Y (n_1571));
  NOR2X1 g37526__4319(.A (n_1566), .B (n_1557), .Y (n_1569));
  OAI21X1 g37494__8428(.A0 (g378), .A1 (n_1552), .B0 (n_1526), .Y
       (n_1568));
  NOR2X1 g37547__5526(.A (n_1566), .B (n_1558), .Y (n_1567));
  NOR4X1 g37872__6783(.A (g1486), .B (g1470), .C (g1504), .D (n_434),
       .Y (n_1565));
  OAI22X1 g37664__3680(.A0 (g321), .A1 (n_1652), .B0 (n_666), .B1
       (n_1662), .Y (n_1580));
  XNOR2X1 g37909__1617(.A (g321), .B (g391), .Y (n_1564));
  OAI21X1 g37911__2802(.A0 (g18), .A1 (n_1563), .B0 (n_1562), .Y
       (n_1573));
  SDFFX1 DFF_230_Q_reg(.CK (CK), .D (n_1548), .SI (n_70), .SE (SE), .Q
       (g342), .QN (n_326));
  SDFFX1 DFF_283_Q_reg(.CK (CK), .D (n_1538), .SI (n_167), .SE (SE), .Q
       (g360), .QN (n_325));
  SDFFX1 DFF_308_Q_reg(.CK (CK), .D (n_1542), .SI (n_22), .SE (SE), .Q
       (g366), .QN (dft_sdo_16));
  SDFFX1 DFF_238_Q_reg(.CK (CK), .D (n_1545), .SI (n_182), .SE (SE), .Q
       (g363), .QN (n_323));
  SDFFX1 DFF_216_Q_reg(.CK (CK), .D (n_1536), .SI (n_176), .SE (SE), .Q
       (g357), .QN (n_322));
  SDFFX1 DFF_499_Q_reg(.CK (CK), .D (n_1540), .SI (n_105), .SE (SE), .Q
       (g339), .QN (n_321));
  INVX1 g37918(.A (n_1562), .Y (n_1575));
  SDFFX1 DFF_490_Q_reg(.CK (CK), .D (n_1530), .SI (g1853), .SE (SE), .Q
       (UNCONNECTED5), .QN (g162));
  NOR2X1 g37511__1705(.A (n_1566), .B (n_1549), .Y (n_1561));
  CLKXOR2X1 g37537__5122(.A (n_1547), .B (n_1544), .Y (n_1560));
  NOR2X1 g37558__8246(.A (n_1570), .B (n_1534), .Y (n_1559));
  AOI22X1 g37560__7098(.A0 (g461), .A1 (n_1556), .B0 (g456), .B1
       (n_1525), .Y (n_1558));
  CLKXOR2X1 g37567__6131(.A (g466), .B (n_1556), .Y (n_1557));
  CLKXOR2X1 g37531__1881(.A (g374), .B (n_1551), .Y (n_1555));
  AND2X1 g37919__5115(.A (g109), .B (g213), .Y (n_1554));
  NAND2X1 g37923__7482(.A (g213), .B (g18), .Y (n_1562));
  NOR2X1 g37548__4733(.A (n_1570), .B (n_1533), .Y (n_1553));
  NOR2X1 g37549__6161(.A (n_401), .B (n_1551), .Y (n_1552));
  NOR2X1 g37565__9315(.A (n_1566), .B (n_1532), .Y (n_1550));
  AOI21X1 g37534__9945(.A0 (g466), .A1 (n_1531), .B0 (g471), .Y
       (n_1549));
  SDFFX1 DFF_478_Q_reg(.CK (CK), .D (g258), .SI (n_73), .SE (SE), .Q
       (UNCONNECTED6), .QN (g321));
  SDFFX1 DFF_430_Q_reg(.CK (CK), .D (n_1523), .SI (n_160), .SE (SE), .Q
       (g481), .QN (n_320));
  SDFFX1 DFF_95_Q_reg(.CK (CK), .D (n_1522), .SI (dft_sdi_5), .SE (SE),
       .Q (g1486), .QN (n_319));
  MX2X1 g37570__2883(.A (g342), .B (n_1546), .S0 (n_1669), .Y (n_1548));
  CLKXOR2X1 g37575__2346(.A (n_1546), .B (n_1541), .Y (n_1547));
  MX2X1 g37564__1666(.A (g363), .B (n_1543), .S0 (n_1669), .Y (n_1545));
  XNOR2X1 g37574__7410(.A (n_1543), .B (n_1537), .Y (n_1544));
  MX2X1 g37573__6417(.A (g366), .B (n_1541), .S0 (n_1669), .Y (n_1542));
  MX2X1 g37568__5477(.A (g339), .B (n_1539), .S0 (n_1669), .Y (n_1540));
  MX2X1 g37571__2398(.A (g360), .B (n_1537), .S0 (n_1669), .Y (n_1538));
  MX2X1 g37569__5107(.A (g357), .B (n_1535), .S0 (n_1669), .Y (n_1536));
  NOR2X1 g37602__6260(.A (g382), .B (n_1527), .Y (n_1534));
  SDFFX1 DFF_447_Q_reg(.CK (CK), .D (n_1505), .SI (n_284), .SE (SE), .Q
       (g521), .QN (n_318));
  SDFFX1 DFF_331_Q_reg(.CK (CK), .D (n_1503), .SI (g1849), .SE (SE), .Q
       (g213), .QN (n_317));
  SDFFX1 DFF_522_Q_reg(.CK (CK), .D (n_1502), .SI (n_166), .SE (SE), .Q
       (g534), .QN (n_316));
  SDFFX1 DFF_368_Q_reg(.CK (CK), .D (n_1511), .SI (n_2), .SE (SE), .Q
       (g448), .QN (n_315));
  SDFFX1 DFF_378_Q_reg(.CK (CK), .D (n_1510), .SI (n_17), .SE (SE), .Q
       (g440), .QN (n_314));
  SDFFX1 DFF_203_Q_reg(.CK (CK), .D (n_1497), .SI (n_103), .SE (SE), .Q
       (g538), .QN (n_313));
  SDFFX1 DFF_492_Q_reg(.CK (CK), .D (n_1492), .SI (n_297), .SE (SE), .Q
       (g431), .QN (n_312));
  SDFFX1 DFF_406_Q_reg(.CK (CK), .D (n_1507), .SI (n_5), .SE (SE), .Q
       (g421), .QN (n_311));
  SDFFX1 DFF_459_Q_reg(.CK (CK), .D (n_1517), .SI (dft_sdi_26), .SE
       (SE), .Q (g506), .QN (n_310));
  SDFFX1 DFF_217_Q_reg(.CK (CK), .D (n_1493), .SI (n_322), .SE (SE), .Q
       (g386), .QN (dft_sdo_11));
  SDFFX1 DFF_3_Q_reg(.CK (CK), .D (n_1512), .SI (g312), .SE (SE), .Q
       (g452), .QN (n_308));
  SDFFX1 DFF_512_Q_reg(.CK (CK), .D (n_1491), .SI (n_89), .SE (SE), .Q
       (g435), .QN (dft_sdo_28));
  SDFFX1 DFF_235_Q_reg(.CK (CK), .D (n_1490), .SI (n_58), .SE (SE), .Q
       (g1432), .QN (dft_sdo_12));
  SDFFX1 DFF_171_Q_reg(.CK (CK), .D (n_1499), .SI (n_42), .SE (SE), .Q
       (g444), .QN (n_305));
  SDFFX1 DFF_210_Q_reg(.CK (CK), .D (n_1494), .SI (n_143), .SE (SE), .Q
       (g530), .QN (n_304));
  SDFFX1 DFF_205_Q_reg(.CK (CK), .D (n_1495), .SI (n_295), .SE (SE), .Q
       (g542), .QN (n_303));
  SDFFX1 DFF_51_Q_reg(.CK (CK), .D (n_1514), .SI (n_161), .SE (SE), .Q
       (g496), .QN (n_302));
  SDFFX1 DFF_419_Q_reg(.CK (CK), .D (n_1506), .SI (n_191), .SE (SE), .Q
       (g406), .QN (n_301));
  SDFFX1 DFF_394_Q_reg(.CK (CK), .D (n_1508), .SI (n_169), .SE (SE), .Q
       (g391), .QN (n_300));
  SDFFX1 DFF_529_Q_reg(.CK (CK), .D (n_1501), .SI (n_156), .SE (SE), .Q
       (g511), .QN (n_299));
  SDFFX1 DFF_475_Q_reg(.CK (CK), .D (n_1518), .SI (g135), .SE (SE), .Q
       (g525), .QN (n_298));
  SDFFX1 DFF_491_Q_reg(.CK (CK), .D (n_1513), .SI (g162), .SE (SE), .Q
       (g411), .QN (n_297));
  SDFFX1 DFF_329_Q_reg(.CK (CK), .D (n_1504), .SI (n_34), .SE (SE), .Q
       (g491), .QN (n_296));
  SDFFX1 DFF_204_Q_reg(.CK (CK), .D (n_1496), .SI (n_313), .SE (SE), .Q
       (g416), .QN (n_295));
  SDFFX1 DFF_221_Q_reg(.CK (CK), .D (n_1519), .SI (n_23), .SE (SE), .Q
       (g501), .QN (n_294));
  SDFFX1 DFF_151_Q_reg(.CK (CK), .D (n_1500), .SI (n_3), .SE (SE), .Q
       (g486), .QN (n_293));
  SDFFX1 DFF_177_Q_reg(.CK (CK), .D (n_1498), .SI (n_85), .SE (SE), .Q
       (g401), .QN (n_292));
  SDFFX1 DFF_379_Q_reg(.CK (CK), .D (n_1509), .SI (n_314), .SE (SE), .Q
       (g476), .QN (n_291));
  SDFFX1 DFF_245_Q_reg(.CK (CK), .D (n_1515), .SI (n_232), .SE (SE), .Q
       (g516), .QN (n_290));
  SDFFX1 DFF_114_Q_reg(.CK (CK), .D (n_1516), .SI (n_52), .SE (SE), .Q
       (g396), .QN (n_289));
  CLKXOR2X1 g37605__4319(.A (g369), .B (n_1528), .Y (n_1533));
  CLKXOR2X1 g37604__8428(.A (g456), .B (n_1524), .Y (n_1532));
  INVX1 g37618(.A (n_1531), .Y (n_1556));
  NAND2X1 g37639__5526(.A (g369), .B (n_1520), .Y (n_1551));
  NOR2X1 g37922__6783(.A (n_1683), .B (n_1736), .Y (n_1530));
  SDFFX1 DFF_206_Q_reg(.CK (CK), .D (n_1489), .SI (n_303), .SE (SE), .Q
       (g560), .QN (n_288));
  SDFFX1 DFF_198_Q_reg(.CK (CK), .D (n_1488), .SI (n_221), .SE (SE), .Q
       (g1346), .QN (dft_sdo_10));
  SDFFX1 DFF_470_Q_reg(.CK (CK), .D (n_1487), .SI (g324), .SE (SE), .Q
       (g1341), .QN (n_286));
  NAND2X1 g37620__3680(.A (g378), .B (n_1528), .Y (n_1529));
  NOR2X1 g37621__1617(.A (n_1526), .B (n_1528), .Y (n_1527));
  NOR2X1 g37623__2802(.A (n_537), .B (n_1524), .Y (n_1525));
  NOR2X1 g37642__1705(.A (n_513), .B (n_1524), .Y (n_1531));
  OAI22X1 g37657__5122(.A0 (n_922), .A1 (n_1662), .B0 (n_650), .B1
       (n_1652), .Y (n_1523));
  OAI22X1 g37659__8246(.A0 (n_710), .A1 (n_1662), .B0 (g309), .B1
       (n_1652), .Y (n_1546));
  OAI22X1 g37662__7098(.A0 (n_622), .A1 (n_1662), .B0 (g333), .B1
       (n_1652), .Y (n_1541));
  SDFFX1 DFF_39_Q_reg(.CK (CK), .D (n_1476), .SI (n_170), .SE (SE), .Q
       (g1543), .QN (dft_sdo_1));
  OAI22X1 g37663__6131(.A0 (g330), .A1 (n_1652), .B0 (n_617), .B1
       (n_1662), .Y (n_1543));
  OAI22X1 g37665__1881(.A0 (g324), .A1 (n_1652), .B0 (n_623), .B1
       (n_1662), .Y (n_1535));
  OAI22X1 g37667__5115(.A0 (n_667), .A1 (n_1662), .B0 (g312), .B1
       (n_1652), .Y (n_1539));
  SDFFX1 DFF_446_Q_reg(.CK (CK), .D (n_1482), .SI (n_18), .SE (SE), .Q
       (g258), .QN (n_284));
  NOR2X1 g37920__7482(.A (n_1683), .B (n_1485), .Y (n_1522));
  CLKINVX2 g37669(.A (n_1528), .Y (n_1520));
  SDFFX1 DFF_249_Q_reg(.CK (CK), .D (n_1479), .SI (n_8), .SE (SE), .Q
       (g1627), .QN (n_283));
  SDFFX1 DFF_133_Q_reg(.CK (CK), .D (n_1473), .SI (n_254), .SE (SE), .Q
       (g281), .QN (n_282));
  OAI22X1 g37668__6161(.A0 (g327), .A1 (n_1652), .B0 (n_698), .B1
       (n_1662), .Y (n_1537));
  SDFFX1 DFF_506_Q_reg(.CK (CK), .D (n_1475), .SI (n_94), .SE (SE), .Q
       (g1351), .QN (n_281));
  MX2X1 g37644__9315(.A (g496), .B (g501), .S0 (n_1662), .Y (n_1519));
  MX2X1 g37622__9945(.A (g530), .B (g525), .S0 (n_1662), .Y (n_1518));
  MX2X1 g37624__2883(.A (g501), .B (g506), .S0 (n_1662), .Y (n_1517));
  MX2X1 g37625__2346(.A (g391), .B (g396), .S0 (n_1662), .Y (n_1516));
  MX2X1 g37626__1666(.A (g511), .B (g516), .S0 (n_1662), .Y (n_1515));
  MX2X1 g37627__7410(.A (g491), .B (g496), .S0 (n_1662), .Y (n_1514));
  MX2X1 g37628__6417(.A (g406), .B (g411), .S0 (n_1662), .Y (n_1513));
  MX2X1 g37629__5477(.A (g421), .B (g452), .S0 (n_1662), .Y (n_1512));
  MX2X1 g37630__2398(.A (g452), .B (g448), .S0 (n_1662), .Y (n_1511));
  MX2X1 g37631__5107(.A (g444), .B (g440), .S0 (n_1662), .Y (n_1510));
  MX2X1 g37632__6260(.A (g516), .B (g476), .S0 (n_1662), .Y (n_1509));
  MX2X1 g37633__4319(.A (g386), .B (g391), .S0 (n_1662), .Y (n_1508));
  MX2X1 g37634__8428(.A (g416), .B (g421), .S0 (n_1662), .Y (n_1507));
  MX2X1 g37635__5526(.A (g401), .B (g406), .S0 (n_1662), .Y (n_1506));
  MX2X1 g37636__6783(.A (g525), .B (g521), .S0 (n_1662), .Y (n_1505));
  MX2X1 g37619__3680(.A (g486), .B (g491), .S0 (n_1662), .Y (n_1504));
  AND2X1 g37942__1617(.A (g109), .B (g1377), .Y (n_1503));
  MX2X1 g37646__2802(.A (g538), .B (g534), .S0 (n_1662), .Y (n_1502));
  MX2X1 g37647__1705(.A (g506), .B (g511), .S0 (n_1662), .Y (n_1501));
  MX2X1 g37648__5122(.A (g481), .B (g486), .S0 (n_1662), .Y (n_1500));
  MX2X1 g37649__8246(.A (g448), .B (g444), .S0 (n_1662), .Y (n_1499));
  MX2X1 g37650__7098(.A (g396), .B (g401), .S0 (n_1662), .Y (n_1498));
  MX2X1 g37651__6131(.A (g542), .B (g538), .S0 (n_1662), .Y (n_1497));
  MX2X1 g37652__1881(.A (g411), .B (g416), .S0 (n_1662), .Y (n_1496));
  MX2X1 g37653__5115(.A (g476), .B (g542), .S0 (n_1662), .Y (n_1495));
  MX2X1 g37654__7482(.A (g534), .B (g530), .S0 (n_1662), .Y (n_1494));
  MX2X1 g37655__4733(.A (g426), .B (g386), .S0 (n_1662), .Y (n_1493));
  MX2X1 g37656__6161(.A (g435), .B (g431), .S0 (n_1662), .Y (n_1492));
  MX2X1 g37645__9315(.A (g440), .B (g435), .S0 (n_1662), .Y (n_1491));
  NOR2X1 g37924__9945(.A (n_1683), .B (n_1481), .Y (n_1490));
  NAND2X1 g37673__2883(.A (n_538), .B (n_1652), .Y (n_1524));
  NAND2X1 g37671__2346(.A (n_1651), .B (n_1652), .Y (n_1528));
  OAI22X1 g37936__1666(.A0 (n_1484), .A1 (n_1586), .B0 (n_1478), .B1
       (n_1631), .Y (n_1489));
  AOI21X1 g37675__7410(.A0 (n_1460), .A1 (n_1471), .B0 (n_1486), .Y
       (n_1488));
  NOR2X1 g37680__6417(.A (n_1486), .B (n_1737), .Y (n_1487));
  XNOR2X1 g37939__5477(.A (n_1484), .B (g1482), .Y (n_1485));
  SDFFX1 DFF_344_Q_reg(.CK (CK), .D (n_1467), .SI (n_12), .SE (SE), .Q
       (g1336), .QN (n_280));
  CLKXOR2X1 g37945__2398(.A (n_1477), .B (g1436), .Y (n_1481));
  SDFFX1 DFF_481_Q_reg(.CK (CK), .D (n_1466), .SI (dft_sdi_27), .SE
       (SE), .Q (g1311), .QN (n_279));
  SDFFX1 DFF_325_Q_reg(.CK (CK), .D (n_1458), .SI (dft_sdi_18), .SE
       (SE), .Q (g1324), .QN (n_278));
  SDFFX1 DFF_458_Q_reg(.CK (CK), .D (n_1463), .SI (n_78), .SE (SE), .Q
       (g1321), .QN (dft_sdo_25));
  SDFFX1 DFF_327_Q_reg(.CK (CK), .D (n_1454), .SI (n_334), .SE (SE), .Q
       (g1377), .QN (n_276));
  CLKINVX2 g37677(.A (n_1662), .Y (n_1652));
  NOR3X1 g37943__5107(.A (n_1047), .B (n_1242), .C (n_1470), .Y
       (n_1480));
  SDFFX1 DFF_448_Q_reg(.CK (CK), .D (n_1462), .SI (n_318), .SE (SE), .Q
       (g1318), .QN (n_275));
  SDFFX1 DFF_195_Q_reg(.CK (CK), .D (n_1461), .SI (g1361), .SE (SE), .Q
       (g1327), .QN (n_274));
  SDFFX1 DFF_146_Q_reg(.CK (CK), .D (n_1457), .SI (n_122), .SE (SE), .Q
       (g1333), .QN (dft_sdo_7));
  SDFFX1 DFF_134_Q_reg(.CK (CK), .D (n_1465), .SI (n_282), .SE (SE), .Q
       (g1308), .QN (n_272));
  SDFFX1 DFF_342_Q_reg(.CK (CK), .D (n_1453), .SI (n_148), .SE (SE), .Q
       (g1314), .QN (n_271));
  SDFFX1 DFF_432_Q_reg(.CK (CK), .D (n_1452), .SI (n_125), .SE (SE), .Q
       (g1330), .QN (n_270));
  MX2X1 g37946__6260(.A (g1627), .B (n_1472), .S0 (n_1631), .Y
       (n_1479));
  OAI21X1 g37960__4319(.A0 (g18), .A1 (n_1478), .B0 (n_1477), .Y
       (n_1482));
  CLKAND2X2 g37679__8428(.A (n_496), .B (n_1468), .Y (n_1662));
  OAI21X1 g37937__5526(.A0 (g1482), .A1 (n_1602), .B0 (n_643), .Y
       (n_1476));
  NOR2X1 g37697__6783(.A (n_1486), .B (n_1469), .Y (n_1475));
  OAI21X1 g37938__1617(.A0 (g174), .A1 (n_1602), .B0 (n_644), .Y
       (n_1473));
  AOI21X1 g37959__2802(.A0 (n_1595), .A1 (g1621), .B0 (n_1472), .Y
       (n_1484));
  NAND3X1 g37685__1705(.A (g1341), .B (n_1443), .C (n_1455), .Y
       (n_1471));
  OAI211X1 g37956__5122(.A0 (g324), .A1 (g396), .B0 (n_1300), .C0
       (n_1357), .Y (n_1470));
  CLKXOR2X1 g37720__8246(.A (g1351), .B (n_1459), .Y (n_1469));
  INVX1 g37970(.A (n_1472), .Y (n_1477));
  NOR4X1 g37682__7098(.A (g841), .B (g853), .C (g857), .D (n_1444), .Y
       (n_1468));
  AND2X1 g37698__6131(.A (n_1451), .B (n_1157), .Y (n_1467));
  SDFFX1 DFF_178_Q_reg(.CK (CK), .D (n_1442), .SI (n_292), .SE (SE), .Q
       (g1857), .QN (n_269));
  MX2X1 g37715__1881(.A (g1771), .B (g1311), .S0 (n_1464), .Y (n_1466));
  MX2X1 g37716__5115(.A (g1766), .B (g1308), .S0 (n_1464), .Y (n_1465));
  MX2X1 g37714__7482(.A (g1786), .B (g1321), .S0 (n_1464), .Y (n_1463));
  MX2X1 g37717__4733(.A (g1781), .B (g1318), .S0 (n_1464), .Y (n_1462));
  MX2X1 g37718__6161(.A (g1796), .B (g1327), .S0 (n_1464), .Y (n_1461));
  NAND2X1 g37721__9315(.A (g1346), .B (n_1459), .Y (n_1460));
  SDFFX1 DFF_102_Q_reg(.CK (CK), .D (n_1439), .SI (n_341), .SE (SE), .Q
       (UNCONNECTED7), .QN (g174));
  SDFFX1 DFF_277_Q_reg(.CK (CK), .D (n_1440), .SI (n_33), .SE (SE), .Q
       (UNCONNECTED8), .QN (g1482));
  MX2X1 g37709__9945(.A (g1791), .B (g1324), .S0 (n_1464), .Y (n_1458));
  MX2X1 g37713__2883(.A (g1806), .B (g1333), .S0 (n_1464), .Y (n_1457));
  SDFFX1 DFF_92_Q_reg(.CK (CK), .D (n_1448), .SI (n_28), .SE (SE), .Q
       (g32), .QN (n_268));
  NOR2X1 g37975__2346(.A (g219), .B (n_1683), .Y (n_1454));
  MX2X1 g37710__1666(.A (g1776), .B (g1314), .S0 (n_1464), .Y (n_1453));
  MX2X1 g37711__7410(.A (g1801), .B (g1330), .S0 (n_1464), .Y (n_1452));
  NOR2X1 g37979__6417(.A (g219), .B (n_1595), .Y (n_1472));
  ADDHX1 g37703__5477(.A (g1336), .B (n_1447), .CO (n_1455), .S
       (n_1451));
  CLKXOR2X1 g37695__2398(.A (n_1449), .B (n_1448), .Y (g11163));
  SDFFX1 DFF_335_Q_reg(.CK (CK), .D (n_1447), .SI (n_102), .SE (SE), .Q
       (g108), .QN (n_267));
  SDFFX1 DFF_420_Q_reg(.CK (CK), .D (n_1435), .SI (n_301), .SE (SE), .Q
       (g1811), .QN (n_266));
  OR2X1 g37706__5107(.A (n_1394), .B (n_1448), .Y (g10801));
  SDFFX1 DFF_467_Q_reg(.CK (CK), .D (g259), .SI (n_74), .SE (SE), .Q
       (UNCONNECTED9), .QN (g324));
  SDFFX1 DFF_125_Q_reg(.CK (CK), .D (n_1430), .SI (n_366), .SE (SE), .Q
       (UNCONNECTED10), .QN (g219));
  NOR4X1 g37935__6260(.A (g237), .B (g231), .C (g225), .D (n_1437), .Y
       (n_1445));
  OR3X1 g37704__4319(.A (g849), .B (g833), .C (n_1436), .Y (n_1444));
  SDFFX1 DFF_73_Q_reg(.CK (CK), .D (n_1433), .SI (n_129), .SE (SE), .Q
       (g563), .QN (n_265));
  OR2X2 g37731__8428(.A (n_1443), .B (n_1438), .Y (n_1459));
  NAND2X1 g37727__5526(.A (g1317), .B (n_1447), .Y (n_1464));
  CLKINVX1 g37712(.A (n_1441), .Y (n_1442));
  SDFFX1 DFF_47_Q_reg(.CK (CK), .D (n_1429), .SI (n_336), .SE (SE), .Q
       (g1436), .QN (n_264));
  AOI222X1 g37719__6783(.A0 (n_506), .A1 (n_928), .B0 (g1857), .B1
       (n_817), .C0 (n_1414), .C1 (n_1427), .Y (n_1441));
  NOR2X1 g37974__3680(.A (n_1683), .B (n_1432), .Y (n_1440));
  NOR2X1 g37976__1617(.A (n_1683), .B (n_1738), .Y (n_1439));
  CLKINVX1 g37735(.A (n_1447), .Y (n_1438));
  SDFFX1 DFF_495_Q_reg(.CK (CK), .D (n_1426), .SI (dft_sdi_28), .SE
       (SE), .Q (g1630), .QN (n_263));
  CLKXOR2X1 g37724__2802(.A (n_500), .B (n_1428), .Y (n_1448));
  NAND4X1 g37971__1705(.A (g1362), .B (g1365), .C (g1368), .D (g1371),
       .Y (n_1437));
  OR4X1 g37728__5122(.A (g837), .B (g829), .C (g861), .D (n_1423), .Y
       (n_1436));
  MX2X1 g37730__8246(.A (g1811), .B (n_1425), .S0 (n_626), .Y (n_1435));
  SDFFX1 DFF_311_Q_reg(.CK (CK), .D (n_1415), .SI (n_184), .SE (SE), .Q
       (g1854), .QN (n_262));
  SDFFX1 DFF_258_Q_reg(.CK (CK), .D (n_1420), .SI (n_95), .SE (SE), .Q
       (g1546), .QN (n_261));
  SDFFX1 DFF_123_Q_reg(.CK (CK), .D (n_1419), .SI (n_65), .SE (SE), .Q
       (g284), .QN (n_260));
  AOI211X1 g37738__7098(.A0 (n_515), .A1 (n_1421), .B0 (n_1384), .C0
       (n_1360), .Y (n_1447));
  OAI22X1 g37988__1881(.A0 (n_1431), .A1 (n_1586), .B0 (n_1411), .B1
       (n_1631), .Y (n_1433));
  CLKXOR2X1 g37992__5115(.A (n_1431), .B (g1478), .Y (n_1432));
  SDFFX1 DFF_193_Q_reg(.CK (CK), .D (n_1416), .SI (n_49), .SE (SE), .Q
       (g259), .QN (n_259));
  NOR2X1 g37997__7482(.A (g1371), .B (n_1683), .Y (n_1430));
  SDFFX1 DFF_120_Q_reg(.CK (CK), .D (n_1408), .SI (n_195), .SE (SE), .Q
       (g1721), .QN (n_258));
  NOR2X1 g37980__4733(.A (n_1683), .B (n_1418), .Y (n_1429));
  CLKXOR2X1 g37737__6161(.A (n_1350), .B (n_1409), .Y (n_1428));
  OAI21X1 g37732__9315(.A0 (n_519), .A1 (n_1344), .B0 (n_1412), .Y
       (n_1427));
  MX2X1 g38002__9945(.A (g1630), .B (n_1413), .S0 (n_1631), .Y
       (n_1426));
  SDFFX1 DFF_67_Q_reg(.CK (CK), .D (n_1403), .SI (n_26), .SE (SE), .Q
       (UNCONNECTED11), .QN (g1371));
  OR4X1 g37741__2883(.A (n_1317), .B (n_1303), .C (n_1424), .D
       (n_1422), .Y (n_1425));
  AOI211X1 g37748__2346(.A0 (g109), .A1 (n_1334), .B0 (n_1363), .C0
       (n_1422), .Y (n_1423));
  NOR4X1 g37750__1666(.A (n_448), .B (n_447), .C (n_558), .D (n_1405),
       .Y (n_1421));
  MX2X1 g37989__7410(.A (g1478), .B (g1546), .S0 (n_1602), .Y (n_1420));
  MX2X1 g37990__6417(.A (g170), .B (g284), .S0 (n_1602), .Y (n_1419));
  CLKXOR2X1 g38000__5477(.A (n_1410), .B (g1440), .Y (n_1418));
  OAI221X1 g37745__2398(.A0 (n_1414), .A1 (n_1319), .B0 (n_1116), .B1
       (n_1400), .C0 (n_1117), .Y (n_1415));
  AOI21X1 g38005__5107(.A0 (n_1595), .A1 (g1624), .B0 (n_1413), .Y
       (n_1431));
  OAI22X1 g37742__6260(.A0 (n_1399), .A1 (n_1402), .B0 (g1690), .B1
       (n_490), .Y (n_1412));
  OAI21X1 g38011__4319(.A0 (g18), .A1 (n_1411), .B0 (n_1410), .Y
       (n_1416));
  CLKXOR2X1 g37749__8428(.A (n_1374), .B (n_1398), .Y (n_1409));
  MX2X1 g37758__5526(.A (n_1407), .B (g1721), .S0 (n_1379), .Y
       (n_1408));
  CLKXOR2X1 g38010__6783(.A (g327), .B (g401), .Y (n_1406));
  INVX1 g38018(.A (n_1410), .Y (n_1413));
  OR3X1 g37767__3680(.A (n_455), .B (n_446), .C (n_1393), .Y (n_1405));
  NAND3X1 g37759__1617(.A (n_1404), .B (n_1378), .C (n_1396), .Y
       (n_1422));
  SDFFX1 DFF_273_Q_reg(.CK (CK), .D (n_1391), .SI (n_215), .SE (SE), .Q
       (g1478), .QN (n_257));
  SDFFX1 DFF_314_Q_reg(.CK (CK), .D (n_1392), .SI (n_147), .SE (SE), .Q
       (g170), .QN (n_256));
  AND2X1 g38021__2802(.A (g109), .B (g225), .Y (n_1403));
  SDFFX1 DFF_168_Q_reg(.CK (CK), .D (n_1401), .SI (g1011), .SE (SE), .Q
       (g33), .QN (n_255));
  NAND2X1 g38023__1705(.A (g225), .B (g18), .Y (n_1410));
  AOI22X1 g37753__5122(.A0 (n_1397), .A1 (n_1401), .B0 (n_1373), .B1
       (n_1376), .Y (n_1402));
  MX2X1 g37766__8246(.A (n_1401), .B (g1806), .S0 (n_1399), .Y
       (n_1400));
  CLKXOR2X1 g37769__7098(.A (n_1397), .B (n_1401), .Y (n_1398));
  INVX1 g37770(.A (n_1396), .Y (n_1407));
  OR2X1 g37774__6131(.A (n_1394), .B (n_1401), .Y (g10455));
  NAND2X1 g37776__1881(.A (g109), .B (n_1401), .Y (n_1396));
  SDFFX1 DFF_65_Q_reg(.CK (CK), .D (g260), .SI (n_124), .SE (SE), .Q
       (UNCONNECTED12), .QN (g327));
  SDFFX1 DFF_132_Q_reg(.CK (CK), .D (n_1381), .SI (n_71), .SE (SE), .Q
       (g225), .QN (n_254));
  SDFFX1 DFF_465_Q_reg(.CK (CK), .D (n_1388), .SI (n_231), .SE (SE), .Q
       (g566), .QN (n_253));
  OAI221X1 g37778__5115(.A0 (g995), .A1 (dft_sdo_26), .B0 (g1250), .B1
       (g1011), .C0 (n_1390), .Y (n_1393));
  SDFFX1 DFF_370_Q_reg(.CK (CK), .D (n_1380), .SI (n_196), .SE (SE), .Q
       (g1727), .QN (n_252));
  SDFFX1 DFF_480_Q_reg(.CK (CK), .D (n_1385), .SI (g321), .SE (SE), .Q
       (UNCONNECTED13), .QN (dft_sdo_26));
  SDFFX1 DFF_503_Q_reg(.CK (CK), .D (n_1377), .SI (n_346), .SE (SE), .Q
       (g1440), .QN (n_251));
  NOR2X1 g38019__7482(.A (n_1683), .B (n_1739), .Y (n_1392));
  NOR2X1 g38020__4733(.A (n_1683), .B (n_1389), .Y (n_1391));
  AOI222X1 g37789__6161(.A0 (n_1361), .A1 (n_1372), .B0 (g995), .B1
       (dft_sdo_26), .C0 (n_1354), .C1 (n_1383), .Y (n_1390));
  SDFFX1 DFF_199_Q_reg(.CK (CK), .D (n_1375), .SI (dft_sdi_11), .SE
       (SE), .Q (g1633), .QN (n_250));
  NAND2X1 g37787__9315(.A (n_960), .B (n_1382), .Y (n_1401));
  SDFFX1 DFF_96_Q_reg(.CK (CK), .D (n_1364), .SI (n_319), .SE (SE), .Q
       (g1730), .QN (n_249));
  SDFFX1 DFF_259_Q_reg(.CK (CK), .D (n_1370), .SI (n_261), .SE (SE), .Q
       (g287), .QN (n_248));
  SDFFX1 DFF_453_Q_reg(.CK (CK), .D (n_1369), .SI (g1393), .SE (SE), .Q
       (g1549), .QN (n_247));
  CLKXOR2X1 g38037__9945(.A (n_1387), .B (g1474), .Y (n_1389));
  OAI22X1 g38034__2883(.A0 (n_1387), .A1 (n_1586), .B0 (n_1359), .B1
       (n_1631), .Y (n_1388));
  SDFFX1 DFF_443_Q_reg(.CK (CK), .D (n_1366), .SI (dft_sdi_25), .SE
       (SE), .Q (g260), .QN (n_246));
  OAI22X1 g37800__1666(.A0 (n_1384), .A1 (n_1383), .B0 (dft_sdo_26),
       .B1 (n_783), .Y (n_1385));
  AOI221X1 g37799__7410(.A0 (n_1296), .A1 (g1567), .B0 (n_1239), .B1
       (g1592), .C0 (n_1362), .Y (n_1382));
  NOR2X1 g38040__6417(.A (g1368), .B (n_1683), .Y (n_1381));
  OAI21X1 g37801__5477(.A0 (n_1379), .A1 (n_1378), .B0 (n_479), .Y
       (n_1380));
  NOR2X1 g38032__2398(.A (n_1683), .B (n_1368), .Y (n_1377));
  SDFFX1 DFF_242_Q_reg(.CK (CK), .D (n_1376), .SI (g330), .SE (SE), .Q
       (g35), .QN (n_245));
  SDFFX1 DFF_530_Q_reg(.CK (CK), .D (n_1356), .SI (n_299), .SE (SE), .Q
       (g1724), .QN (n_244));
  MX2X1 g38051__5107(.A (g1633), .B (n_1365), .S0 (n_1631), .Y
       (n_1375));
  SDFFX1 DFF_163_Q_reg(.CK (CK), .D (n_1353), .SI (n_243), .SE (SE), .Q
       (UNCONNECTED14), .QN (g1368));
  CLKXOR2X1 g37814__6260(.A (n_1373), .B (n_1376), .Y (n_1374));
  CLKINVX2 g37825(.A (n_1383), .Y (n_1372));
  OR2X1 g37818__4319(.A (n_1394), .B (n_1376), .Y (g10459));
  OAI21X1 g38031__8428(.A0 (g127), .A1 (n_1602), .B0 (n_641), .Y
       (n_1370));
  MX2X1 g38036__5526(.A (g1474), .B (g1549), .S0 (n_1602), .Y (n_1369));
  CLKXOR2X1 g38046__6783(.A (n_1358), .B (g1444), .Y (n_1368));
  AOI21X1 g38067__3680(.A0 (n_1595), .A1 (g1627), .B0 (n_1365), .Y
       (n_1387));
  MX2X1 g37813__1617(.A (n_1363), .B (g1730), .S0 (n_1379), .Y
       (n_1364));
  NAND2X1 g37830__2802(.A (n_958), .B (n_1355), .Y (n_1362));
  SDFFX1 DFF_161_Q_reg(.CK (CK), .D (n_1351), .SI (n_117), .SE (SE), .Q
       (g105), .QN (n_243));
  AOI22X1 g37815__1705(.A0 (g109), .A1 (n_1290), .B0 (g108), .B1
       (n_1363), .Y (n_1449));
  NAND2X1 g37820__5122(.A (g109), .B (n_1376), .Y (n_1378));
  MX2X1 g37833__8246(.A (n_909), .B (n_1361), .S0 (n_1360), .Y
       (n_1383));
  OAI21X1 g38068__7098(.A0 (g18), .A1 (n_1359), .B0 (n_1358), .Y
       (n_1366));
  CLKXOR2X1 g38065__6131(.A (g330), .B (g406), .Y (n_1357));
  SDFFX1 DFF_228_Q_reg(.CK (CK), .D (n_1373), .SI (n_159), .SE (SE), .Q
       (g36), .QN (n_242));
  INVX1 g38078(.A (n_1358), .Y (n_1365));
  OAI21X1 g37845__1881(.A0 (n_1379), .A1 (n_1404), .B0 (n_475), .Y
       (n_1356));
  AOI221X1 g37842__5115(.A0 (g898), .A1 (n_1347), .B0 (g922), .B1
       (n_1051), .C0 (n_1346), .Y (n_1355));
  INVX1 g37854(.A (n_1361), .Y (n_1354));
  NAND4X1 g37840__7482(.A (n_1066), .B (n_1345), .C (n_962), .D
       (n_1348), .Y (n_1376));
  AND2X1 g38081__4733(.A (g109), .B (g231), .Y (n_1353));
  SDFFX1 DFF_508_Q_reg(.CK (CK), .D (n_1340), .SI (n_281), .SE (SE), .Q
       (UNCONNECTED15), .QN (g127));
  NAND2X1 g38088__6161(.A (g231), .B (g18), .Y (n_1358));
  SDFFX1 DFF_172_Q_reg(.CK (CK), .D (n_1341), .SI (n_305), .SE (SE), .Q
       (g1474), .QN (n_241));
  SDFFX1 DFF_384_Q_reg(.CK (CK), .D (n_1397), .SI (n_134), .SE (SE), .Q
       (g34), .QN (n_240));
  SDFFX1 DFF_423_Q_reg(.CK (CK), .D (n_1342), .SI (n_266), .SE (SE), .Q
       (g1654), .QN (n_239));
  CLKINVX2 g37841(.A (n_1424), .Y (n_1363));
  CLKXOR2X1 g37858__9315(.A (g1027), .B (n_1343), .Y (n_1361));
  OR2X1 g37838__9945(.A (n_1394), .B (n_1373), .Y (g10461));
  MX2X1 g37855__2883(.A (g105), .B (n_1339), .S0 (n_1631), .Y (n_1351));
  NAND2X1 g37848__2346(.A (g109), .B (n_1373), .Y (n_1424));
  CLKXOR2X1 g37847__1666(.A (n_1328), .B (n_1277), .Y (n_1350));
  OR2X1 g37860__7410(.A (n_1394), .B (n_1397), .Y (g10457));
  SDFFX1 DFF_239_Q_reg(.CK (CK), .D (g261), .SI (n_323), .SE (SE), .Q
       (UNCONNECTED16), .QN (g330));
  SDFFX1 DFF_185_Q_reg(.CK (CK), .D (n_1318), .SI (n_157), .SE (SE), .Q
       (g231), .QN (n_238));
  AOI221X1 g37874__6417(.A0 (n_1265), .A1 (g269), .B0 (g904), .B1
       (n_1347), .C0 (n_1330), .Y (n_1348));
  NAND3X1 g37867__5477(.A (n_1309), .B (n_1345), .C (n_1327), .Y
       (n_1346));
  SDFFX1 DFF_524_Q_reg(.CK (CK), .D (n_1325), .SI (n_97), .SE (SE), .Q
       (g569), .QN (n_237));
  NAND2X1 g37865__2398(.A (g109), .B (n_1397), .Y (n_1404));
  NOR2X1 g37837__5107(.A (n_1399), .B (n_1337), .Y (n_1344));
  NAND2X1 g37859__6260(.A (n_996), .B (n_1335), .Y (n_1373));
  NAND2X1 g37878__4319(.A (g1032), .B (n_1329), .Y (n_1343));
  SDFFX1 DFF_36_Q_reg(.CK (CK), .D (n_1316), .SI (n_364), .SE (SE), .Q
       (g1444), .QN (n_236));
  MX2X1 g38083__8428(.A (n_1315), .B (g1654), .S0 (n_1251), .Y
       (n_1342));
  NOR2X1 g38082__5526(.A (n_1683), .B (n_1323), .Y (n_1341));
  NOR2X1 g38080__6783(.A (n_1683), .B (n_1740), .Y (n_1340));
  OR2X1 g37876__3680(.A (n_881), .B (n_1338), .Y (n_1339));
  SDFFX1 DFF_22_Q_reg(.CK (CK), .D (n_1336), .SI (n_79), .SE (SE), .Q
       (g39), .QN (n_235));
  SDFFX1 DFF_251_Q_reg(.CK (CK), .D (n_1313), .SI (n_104), .SE (SE), .Q
       (g290), .QN (n_234));
  SDFFX1 DFF_404_Q_reg(.CK (CK), .D (n_1312), .SI (n_126), .SE (SE), .Q
       (g1636), .QN (dft_sdo_22));
  NAND3X1 g37888__1617(.A (n_1345), .B (n_957), .C (n_1314), .Y
       (n_1397));
  AOI22X1 g37856__2802(.A0 (n_1332), .A1 (n_1331), .B0 (n_1333), .B1
       (n_1336), .Y (n_1337));
  AOI221X1 g37871__1705(.A0 (g1203), .A1 (n_1320), .B0 (g8), .B1
       (n_1287), .C0 (n_1311), .Y (n_1335));
  OR4X1 g37882__5122(.A (n_1333), .B (n_1332), .C (n_1331), .D
       (n_1336), .Y (n_1334));
  INVX1 g37895(.A (n_1321), .Y (n_1330));
  INVX1 g37889(.A (n_1338), .Y (n_1329));
  XNOR2X1 g37887__8246(.A (n_1333), .B (n_1336), .Y (n_1328));
  AOI221X1 g37897__7098(.A0 (n_1087), .A1 (g971), .B0 (n_1222), .B1
       (g33), .C0 (n_1310), .Y (n_1327));
  OAI22X1 g38116__1881(.A0 (n_1322), .A1 (n_1586), .B0 (n_1299), .B1
       (n_1631), .Y (n_1325));
  OR2X1 g37890__5115(.A (n_1394), .B (n_1336), .Y (g10377));
  XNOR2X1 g38120__7482(.A (n_1322), .B (g1470), .Y (n_1323));
  SDFFX1 DFF_244_Q_reg(.CK (CK), .D (n_1306), .SI (n_245), .SE (SE), .Q
       (g261), .QN (n_232));
  AOI221X1 g37896__4733(.A0 (n_1286), .A1 (g293), .B0 (g1200), .B1
       (n_1320), .C0 (n_1305), .Y (n_1321));
  OAI21X1 g37901__6161(.A0 (n_745), .A1 (n_1304), .B0 (g1854), .Y
       (n_1319));
  NOR2X1 g38129__9315(.A (g1365), .B (n_1683), .Y (n_1318));
  SDFFX1 DFF_463_Q_reg(.CK (CK), .D (n_1301), .SI (n_217), .SE (SE), .Q
       (g1552), .QN (n_231));
  NOR2X1 g37894__9945(.A (n_1317), .B (n_1336), .Y (n_1338));
  NOR2X1 g38095__2883(.A (n_1683), .B (n_1308), .Y (n_1316));
  NOR2X1 g38128__2346(.A (g1718), .B (n_1322), .Y (n_1315));
  AOI221X1 g37910__1666(.A0 (n_1294), .A1 (g1341), .B0 (g1173), .B1
       (n_1284), .C0 (n_1292), .Y (n_1314));
  SDFFX1 DFF_321_Q_reg(.CK (CK), .D (n_1289), .SI (n_227), .SE (SE), .Q
       (g1733), .QN (n_230));
  MX2X1 g38117__7410(.A (g131), .B (g290), .S0 (n_1602), .Y (n_1313));
  MX2X1 g38147__6417(.A (g1636), .B (n_1302), .S0 (n_1631), .Y
       (n_1312));
  SDFFX1 DFF_142_Q_reg(.CK (CK), .D (n_1280), .SI (n_116), .SE (SE), .Q
       (UNCONNECTED17), .QN (g1365));
  NAND2X1 g37898__5477(.A (n_1057), .B (n_1297), .Y (n_1311));
  OAI211X1 g37907__2398(.A0 (n_1190), .A1 (n_395), .B0 (n_1077), .C0
       (n_1288), .Y (n_1310));
  NAND3X1 g37912__5107(.A (n_1309), .B (n_1059), .C (n_1285), .Y
       (n_1336));
  CLKXOR2X1 g38148__6260(.A (n_1298), .B (g1448), .Y (n_1308));
  INVX1 g37917(.A (n_1295), .Y (n_1305));
  OAI211X1 g37934__4319(.A0 (n_1281), .A1 (n_1303), .B0 (n_702), .C0
       (n_1282), .Y (n_1304));
  AOI21X1 g38174__8428(.A0 (n_1595), .A1 (g1630), .B0 (n_1302), .Y
       (n_1322));
  OAI21X1 g38118__5526(.A0 (g1470), .A1 (n_1602), .B0 (n_640), .Y
       (n_1301));
  CLKXOR2X1 g38166__6783(.A (g333), .B (g411), .Y (n_1300));
  OAI21X1 g38173__3680(.A0 (g18), .A1 (n_1299), .B0 (n_1298), .Y
       (n_1306));
  AOI221X1 g37908__1617(.A0 (n_1296), .A1 (g1577), .B0 (n_1293), .B1
       (g1730), .C0 (n_1273), .Y (n_1297));
  AOI221X1 g37921__2802(.A0 (n_1294), .A1 (g1346), .B0 (n_1293), .B1
       (g1727), .C0 (n_1275), .Y (n_1295));
  OAI211X1 g37926__1705(.A0 (n_1034), .A1 (n_1291), .B0 (n_1095), .C0
       (n_1276), .Y (n_1292));
  INVX1 g37944(.A (n_1283), .Y (n_1290));
  MX2X1 g37947__5122(.A (n_1303), .B (g1733), .S0 (n_1379), .Y
       (n_1289));
  SDFFX1 DFF_444_Q_reg(.CK (CK), .D (n_1267), .SI (n_246), .SE (SE), .Q
       (g131), .QN (n_229));
  AOI221X1 g37933__8246(.A0 (n_1287), .A1 (g123), .B0 (n_1286), .B1
       (g287), .C0 (n_1271), .Y (n_1288));
  AOI221X1 g37940__7098(.A0 (n_1171), .A1 (g1333), .B0 (g1188), .B1
       (n_1284), .C0 (n_1270), .Y (n_1285));
  INVX1 g38176(.A (n_1298), .Y (n_1302));
  AOI222X1 g37948__6131(.A0 (g2648), .A1 (n_1333), .B0 (n_918), .B1
       (n_1332), .C0 (n_388), .C1 (n_1331), .Y (n_1283));
  NAND2X1 g37950__1881(.A (n_1281), .B (n_1303), .Y (n_1282));
  AND2X1 g38183__5115(.A (g109), .B (g237), .Y (n_1280));
  SDFFX1 DFF_350_Q_reg(.CK (CK), .D (n_1332), .SI (n_145), .SE (SE), .Q
       (g37), .QN (n_228));
  NAND2X1 g38198__7482(.A (g237), .B (g18), .Y (n_1298));
  NOR2X1 g37972__4733(.A (n_1278), .B (n_1268), .Y (n_1279));
  CLKXOR2X1 g37958__6161(.A (n_1332), .B (n_1331), .Y (n_1277));
  AND3X2 g37957__9315(.A (n_993), .B (n_1162), .C (n_1274), .Y
       (n_1276));
  SDFFX1 DFF_319_Q_reg(.CK (CK), .D (n_1333), .SI (n_113), .SE (SE), .Q
       (g40), .QN (n_227));
  NAND4X1 g37925__9945(.A (n_995), .B (n_1069), .C (n_1038), .D
       (n_1274), .Y (n_1275));
  NAND4X1 g37927__2883(.A (n_961), .B (n_999), .C (n_1168), .D
       (n_1274), .Y (n_1273));
  SDFFX1 DFF_175_Q_reg(.CK (CK), .D (g262), .SI (n_121), .SE (SE), .Q
       (UNCONNECTED18), .QN (g333));
  SDFFX1 DFF_98_Q_reg(.CK (CK), .D (n_1263), .SI (g1504), .SE (SE), .Q
       (UNCONNECTED19), .QN (g1470));
  OR2X1 g37973__2346(.A (n_1394), .B (n_1332), .Y (g10463));
  NAND2X1 g37949__1666(.A (n_1049), .B (n_1274), .Y (n_1271));
  NAND2X1 g37955__7410(.A (n_994), .B (n_1266), .Y (n_1270));
  SDFFX1 DFF_166_Q_reg(.CK (CK), .D (n_1260), .SI (dft_sdi_9), .SE
       (SE), .Q (g572), .QN (n_226));
  SDFFX1 DFF_303_Q_reg(.CK (CK), .D (n_1258), .SI (n_187), .SE (SE), .Q
       (g237), .QN (n_225));
  OR2X1 g37968__6417(.A (n_1683), .B (n_1332), .Y (n_1303));
  OR2X1 g37963__5477(.A (n_1394), .B (n_1333), .Y (g10379));
  INVX1 g37986(.A (n_1332), .Y (n_1268));
  NOR2X1 g38178__2398(.A (n_1683), .B (n_1741), .Y (n_1267));
  SDFFX1 DFF_116_Q_reg(.CK (CK), .D (n_1331), .SI (n_56), .SE (SE), .Q
       (g38), .QN (n_224));
  SDFFX1 DFF_285_Q_reg(.CK (CK), .D (n_1252), .SI (g192), .SE (SE), .Q
       (g1657), .QN (n_223));
  AOI221X1 g37977__5107(.A0 (n_1265), .A1 (g281), .B0 (g916), .B1
       (n_1347), .C0 (n_1257), .Y (n_1266));
  OR3X1 g37978__6260(.A (n_1320), .B (n_1294), .C (n_1264), .Y
       (n_1274));
  SDFFX1 DFF_360_Q_reg(.CK (CK), .D (n_1250), .SI (n_202), .SE (SE), .Q
       (g636), .QN (n_222));
  SDFFX1 DFF_197_Q_reg(.CK (CK), .D (n_1249), .SI (n_133), .SE (SE), .Q
       (g293), .QN (n_221));
  NAND4X1 g37993__4319(.A (n_955), .B (n_1092), .C (n_1205), .D
       (n_1264), .Y (n_1332));
  NOR2X1 g38179__8428(.A (n_1683), .B (n_1254), .Y (n_1263));
  NAND2X1 g37985__6783(.A (n_1088), .B (n_1256), .Y (n_1333));
  SDFFX1 DFF_222_Q_reg(.CK (CK), .D (n_1247), .SI (n_294), .SE (SE), .Q
       (g262), .QN (n_220));
  OR2X1 g37994__3680(.A (n_1394), .B (n_1331), .Y (g10465));
  SDFFX1 DFF_191_Q_reg(.CK (CK), .D (n_1245), .SI (n_343), .SE (SE), .Q
       (g627), .QN (n_219));
  OAI221X1 g38215__1617(.A0 (n_1253), .A1 (n_1149), .B0 (n_1244), .B1
       (n_1631), .C0 (n_1259), .Y (n_1260));
  NOR2X1 g38304__2802(.A (g1362), .B (n_1683), .Y (n_1258));
  SDFFX1 DFF_514_Q_reg(.CK (CK), .D (n_1243), .SI (dft_sdi_29), .SE
       (SE), .Q (g1555), .QN (n_218));
  OAI21X1 g37999__1705(.A0 (n_1294), .A1 (n_1255), .B0 (n_959), .Y
       (n_1257));
  AOI21X1 g38001__5122(.A0 (n_1296), .A1 (g1589), .B0 (n_1246), .Y
       (n_1256));
  OR3X1 g38003__8246(.A (n_1287), .B (n_1204), .C (n_1255), .Y
       (n_1264));
  XNOR2X1 g38274__7098(.A (n_1253), .B (g1466), .Y (n_1254));
  OAI211X1 g38216__6131(.A0 (n_1251), .A1 (n_1253), .B0 (n_504), .C0
       (n_1119), .Y (n_1252));
  SDFFX1 DFF_461_Q_reg(.CK (CK), .D (n_1241), .SI (n_310), .SE (SE), .Q
       (g1909), .QN (n_217));
  NAND3X1 g38012__1881(.A (n_1003), .B (n_1255), .C (n_1240), .Y
       (n_1331));
  OAI222X1 g38204__5115(.A0 (n_595), .A1 (n_1099), .B0 (n_1113), .B1
       (n_1238), .C0 (g622), .C1 (n_1042), .Y (n_1250));
  OAI21X1 g38272__7482(.A0 (g135), .A1 (n_1602), .B0 (n_645), .Y
       (n_1249));
  SDFFX1 DFF_88_Q_reg(.CK (CK), .D (n_1226), .SI (n_48), .SE (SE), .Q
       (UNCONNECTED20), .QN (g1362));
  SDFFX1 DFF_354_Q_reg(.CK (CK), .D (n_1227), .SI (n_139), .SE (SE), .Q
       (g1891), .QN (n_216));
  SDFFX1 DFF_271_Q_reg(.CK (CK), .D (n_1229), .SI (dft_sdi_15), .SE
       (SE), .Q (g1945), .QN (n_215));
  SDFFX1 DFF_44_Q_reg(.CK (CK), .D (n_1235), .SI (n_186), .SE (SE), .Q
       (g1927), .QN (n_214));
  SDFFX1 DFF_1_Q_reg(.CK (CK), .D (n_1232), .SI (scan_in), .SE (SE), .Q
       (g1882), .QN (n_213));
  SDFFX1 DFF_300_Q_reg(.CK (CK), .D (n_1225), .SI (n_152), .SE (SE), .Q
       (g1918), .QN (n_212));
  SDFFX1 DFF_212_Q_reg(.CK (CK), .D (n_1223), .SI (n_190), .SE (SE), .Q
       (g1936), .QN (n_211));
  SDFFX1 DFF_449_Q_reg(.CK (CK), .D (n_1224), .SI (n_275), .SE (SE), .Q
       (g1872), .QN (n_210));
  SDFFX1 DFF_333_Q_reg(.CK (CK), .D (n_1228), .SI (n_96), .SE (SE), .Q
       (g1900), .QN (n_209));
  OAI211X1 g38009__4733(.A0 (n_1294), .A1 (n_1234), .B0 (n_1056), .C0
       (n_1000), .Y (n_1246));
  NOR2X1 g38312__6161(.A (g635), .B (n_1209), .Y (n_1245));
  OAI21X1 g38371__9315(.A0 (g18), .A1 (n_1244), .B0 (n_1237), .Y
       (n_1247));
  OAI21X1 g38271__9945(.A0 (g1466), .A1 (n_1602), .B0 (n_637), .Y
       (n_1243));
  OAI211X1 g38022__2883(.A0 (n_887), .A1 (n_858), .B0 (n_893), .C0
       (n_1233), .Y (n_1255));
  XNOR2X1 g38359__2346(.A (g309), .B (g416), .Y (n_1242));
  AOI21X1 g38373__1666(.A0 (n_1595), .A1 (g1633), .B0 (n_1236), .Y
       (n_1253));
  INVX1 g38105(.A (n_1230), .Y (n_1241));
  AOI221X1 g38145__7410(.A0 (n_1239), .A1 (g1607), .B0 (g1185), .B1
       (n_1284), .C0 (n_1221), .Y (n_1240));
  SDFFX1 DFF_362_Q_reg(.CK (CK), .D (n_1217), .SI (n_192), .SE (SE), .Q
       (g605), .QN (n_208));
  SDFFX1 DFF_135_Q_reg(.CK (CK), .D (n_1214), .SI (n_272), .SE (SE), .Q
       (g611), .QN (n_207));
  SDFFX1 DFF_157_Q_reg(.CK (CK), .D (n_1219), .SI (n_151), .SE (SE), .Q
       (UNCONNECTED21), .QN (g635));
  OAI21X1 g38282__6417(.A0 (n_1220), .A1 (n_1048), .B0 (g636), .Y
       (n_1238));
  CLKINVX1 g38381(.A (n_1236), .Y (n_1237));
  SDFFX1 DFF_474_Q_reg(.CK (CK), .D (n_1215), .SI (n_369), .SE (SE), .Q
       (UNCONNECTED22), .QN (g135));
  SDFFX1 DFF_455_Q_reg(.CK (CK), .D (n_1216), .SI (n_382), .SE (SE), .Q
       (g1834), .QN (n_206));
  OAI211X1 g38109__5477(.A0 (n_717), .A1 (n_1213), .B0 (n_1186), .C0
       (n_1231), .Y (n_1235));
  INVX1 g38045(.A (n_1233), .Y (n_1234));
  OAI211X1 g38143__2398(.A0 (n_938), .A1 (n_1203), .B0 (n_1189), .C0
       (n_1231), .Y (n_1232));
  AOI221X1 g38107__5107(.A0 (n_1019), .A1 (n_1118), .B0 (g1909), .B1
       (n_1187), .C0 (n_1151), .Y (n_1230));
  OAI211X1 g38108__6260(.A0 (n_800), .A1 (n_1218), .B0 (n_1181), .C0
       (n_1231), .Y (n_1229));
  OAI211X1 g38137__4319(.A0 (n_932), .A1 (n_1208), .B0 (n_1179), .C0
       (n_1231), .Y (n_1228));
  OAI211X1 g38110__8428(.A0 (n_469), .A1 (n_1210), .B0 (n_1183), .C0
       (n_1231), .Y (n_1227));
  NOR2X1 g38395__5526(.A (g243), .B (n_1683), .Y (n_1226));
  SDFFX1 DFF_6_Q_reg(.CK (CK), .D (n_1195), .SI (n_342), .SE (SE), .Q
       (g713), .QN (n_205));
  NOR2X1 g38398__6783(.A (g243), .B (n_1595), .Y (n_1236));
  SDFFX1 DFF_395_Q_reg(.CK (CK), .D (n_1192), .SI (n_300), .SE (SE), .Q
       (g658), .QN (n_204));
  OAI211X1 g38146__3680(.A0 (n_935), .A1 (n_1206), .B0 (n_1174), .C0
       (n_1231), .Y (n_1225));
  OAI211X1 g38149__1617(.A0 (n_470), .A1 (n_1202), .B0 (n_1170), .C0
       (n_1231), .Y (n_1224));
  OAI211X1 g38144__2802(.A0 (n_937), .A1 (n_1207), .B0 (n_1176), .C0
       (n_1231), .Y (n_1223));
  SDFFX1 DFF_11_Q_reg(.CK (CK), .D (n_1197), .SI (n_155), .SE (SE), .Q
       (g695), .QN (n_203));
  SDFFX1 DFF_359_Q_reg(.CK (CK), .D (n_1200), .SI (n_188), .SE (SE), .Q
       (g731), .QN (n_202));
  SDFFX1 DFF_57_Q_reg(.CK (CK), .D (n_1196), .SI (n_40), .SE (SE), .Q
       (g704), .QN (dft_sdo_2));
  SDFFX1 DFF_316_Q_reg(.CK (CK), .D (n_1194), .SI (n_21), .SE (SE), .Q
       (g686), .QN (n_200));
  SDFFX1 DFF_450_Q_reg(.CK (CK), .D (n_1198), .SI (n_210), .SE (SE), .Q
       (g677), .QN (n_199));
  SDFFX1 DFF_286_Q_reg(.CK (CK), .D (n_1201), .SI (n_223), .SE (SE), .Q
       (g722), .QN (n_198));
  SDFFX1 DFF_381_Q_reg(.CK (CK), .D (n_1193), .SI (n_32), .SE (SE), .Q
       (g668), .QN (n_197));
  SDFFX1 DFF_369_Q_reg(.CK (CK), .D (n_1177), .SI (n_315), .SE (SE), .Q
       (g1828), .QN (n_196));
  NOR4X1 g38052__1705(.A (n_1222), .B (n_1296), .C (n_1347), .D
       (n_1191), .Y (n_1233));
  SDFFX1 DFF_183_Q_reg(.CK (CK), .D (g254), .SI (n_158), .SE (SE), .Q
       (UNCONNECTED23), .QN (g309));
  SDFFX1 DFF_119_Q_reg(.CK (CK), .D (n_1167), .SI (n_20), .SE (SE), .Q
       (g1227), .QN (n_195));
  SDFFX1 DFF_139_Q_reg(.CK (CK), .D (n_1160), .SI (n_69), .SE (SE), .Q
       (UNCONNECTED24), .QN (g1466));
  SDFFX1 DFF_28_Q_reg(.CK (CK), .D (n_1159), .SI (n_37), .SE (SE), .Q
       (g1231), .QN (n_194));
  SDFFX1 DFF_297_Q_reg(.CK (CK), .D (n_1161), .SI (n_180), .SE (SE), .Q
       (g1814), .QN (n_193));
  SDFFX1 DFF_361_Q_reg(.CK (CK), .D (n_1164), .SI (n_222), .SE (SE), .Q
       (g1218), .QN (n_192));
  SDFFX1 DFF_418_Q_reg(.CK (CK), .D (n_1158), .SI (n_338), .SE (SE), .Q
       (g1223), .QN (n_191));
  NAND2X1 g38200__5122(.A (n_1058), .B (n_1172), .Y (n_1221));
  SDFFX1 DFF_33_Q_reg(.CK (CK), .D (n_1153), .SI (n_106), .SE (SE), .Q
       (UNCONNECTED25), .QN (g243));
  CLKINVX1 g38380(.A (n_1219), .Y (n_1220));
  SDFFX1 DFF_211_Q_reg(.CK (CK), .D (n_1150), .SI (n_304), .SE (SE), .Q
       (g575), .QN (n_190));
  AOI21X1 g38201__8246(.A0 (n_1180), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1218));
  AND2X1 g38090__7098(.A (n_1165), .B (g18), .Y (n_1217));
  AOI21X1 g38167__6131(.A0 (n_832), .A1 (n_1155), .B0 (n_1595), .Y
       (n_1216));
  NOR2X1 g38394__1881(.A (n_1683), .B (n_1742), .Y (n_1215));
  AOI21X1 g38084__5115(.A0 (n_869), .A1 (n_1154), .B0 (n_1595), .Y
       (n_1214));
  AOI21X1 g38202__7482(.A0 (n_1185), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1213));
  AOI21X1 g38203__4733(.A0 (n_1182), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1210));
  NOR2X1 g38397__6161(.A (g632), .B (n_1209), .Y (n_1219));
  AOI21X1 g38224__9315(.A0 (n_1178), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1208));
  AOI21X1 g38227__9945(.A0 (n_1175), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1207));
  AOI21X1 g38229__2883(.A0 (n_1173), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1206));
  AOI221X1 g38236__2346(.A0 (n_1037), .A1 (g962), .B0 (g16), .B1
       (n_1204), .C0 (n_1148), .Y (n_1205));
  AOI21X1 g38226__1666(.A0 (n_1188), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1203));
  AOI21X1 g38260__7410(.A0 (n_1169), .A1 (n_1212), .B0 (n_1211), .Y
       (n_1202));
  SDFFX1 DFF_45_Q_reg(.CK (CK), .D (n_1120), .SI (n_214), .SE (SE), .Q
       (g1660), .QN (n_189));
  SDFFX1 DFF_358_Q_reg(.CK (CK), .D (n_1128), .SI (n_136), .SE (SE), .Q
       (g591), .QN (n_188));
  SDFFX1 DFF_302_Q_reg(.CK (CK), .D (n_1125), .SI (n_140), .SE (SE), .Q
       (g1822), .QN (n_187));
  OAI211X1 g38063__6417(.A0 (n_1046), .A1 (n_1108), .B0 (n_1129), .C0
       (n_1199), .Y (n_1201));
  OAI211X1 g38048__5477(.A0 (n_776), .A1 (n_1140), .B0 (n_1136), .C0
       (n_1199), .Y (n_1200));
  OAI211X1 g38049__2398(.A0 (n_405), .A1 (n_1143), .B0 (n_1134), .C0
       (n_1199), .Y (n_1198));
  OAI211X1 g38050__5107(.A0 (n_548), .A1 (n_1144), .B0 (n_1131), .C0
       (n_1199), .Y (n_1197));
  OAI211X1 g38061__6260(.A0 (n_649), .A1 (n_1086), .B0 (n_1145), .C0
       (n_1199), .Y (n_1196));
  OAI211X1 g38047__4319(.A0 (n_688), .A1 (n_1106), .B0 (n_1132), .C0
       (n_1199), .Y (n_1195));
  OAI211X1 g38064__8428(.A0 (n_1045), .A1 (n_1104), .B0 (n_1139), .C0
       (n_1199), .Y (n_1194));
  OAI211X1 g38066__5526(.A0 (n_1043), .A1 (n_1110), .B0 (n_1137), .C0
       (n_1199), .Y (n_1193));
  OAI211X1 g38111__6783(.A0 (n_904), .A1 (n_1080), .B0 (n_1126), .C0
       (n_1199), .Y (n_1192));
  NAND4X1 g38121__3680(.A (n_949), .B (n_1190), .C (n_890), .D
       (n_1127), .Y (n_1191));
  SDFFX1 DFF_43_Q_reg(.CK (CK), .D (n_1114), .SI (n_83), .SE (SE), .Q
       (g622), .QN (n_186));
  OR3X1 g38257__1617(.A (g1882), .B (n_1188), .C (n_1184), .Y (n_1189));
  OAI21X1 g38207__2802(.A0 (n_970), .A1 (n_1115), .B0 (n_1156), .Y
       (n_1187));
  OR3X1 g38208__1705(.A (g1927), .B (n_1185), .C (n_1184), .Y (n_1186));
  OR3X1 g38209__5122(.A (g1891), .B (n_1182), .C (n_1184), .Y (n_1183));
  OR3X1 g38210__8246(.A (g1945), .B (n_1180), .C (n_1184), .Y (n_1181));
  OR3X1 g38256__7098(.A (g1900), .B (n_1178), .C (n_1184), .Y (n_1179));
  AND2X1 g38181__6131(.A (n_1152), .B (g18), .Y (n_1177));
  OR3X1 g38258__1881(.A (g1936), .B (n_1175), .C (n_1184), .Y (n_1176));
  OR3X1 g38266__5115(.A (g1918), .B (n_1173), .C (n_1184), .Y (n_1174));
  AOI221X1 g38270__7482(.A0 (n_1171), .A1 (g1330), .B0 (n_1286), .B1
       (g302), .C0 (n_1121), .Y (n_1172));
  OR3X1 g38303__4733(.A (g1872), .B (n_1169), .C (n_1184), .Y (n_1170));
  AOI221X1 g38308__6161(.A0 (n_1222), .A1 (g36), .B0 (g17), .B1
       (n_1204), .C0 (n_1122), .Y (n_1168));
  AOI21X1 g38233__9315(.A0 (n_695), .A1 (n_868), .B0 (n_1163), .Y
       (n_1167));
  SDFFX1 DFF_246_Q_reg(.CK (CK), .D (n_1111), .SI (n_290), .SE (SE), .Q
       (g254), .QN (n_185));
  SDFFX1 DFF_117_Q_reg(.CK (CK), .D (n_1091), .SI (n_224), .SE (SE), .Q
       (UNCONNECTED26), .QN (g632));
  CLKXOR2X1 g38136__2883(.A (g605), .B (n_1100), .Y (n_1165));
  NOR2X1 g38393__2346(.A (n_1163), .B (n_739), .Y (n_1164));
  AOI21X1 g38230__1666(.A0 (n_1293), .A1 (g1724), .B0 (n_1123), .Y
       (n_1162));
  AND2X1 g38232__7410(.A (n_1124), .B (g18), .Y (n_1161));
  SDFFX1 DFF_310_Q_reg(.CK (CK), .D (n_1094), .SI (n_4), .SE (SE), .Q
       (g599), .QN (n_184));
  SDFFX1 DFF_252_Q_reg(.CK (CK), .D (n_1090), .SI (n_234), .SE (SE), .Q
       (g1850), .QN (n_183));
  NOR2X1 g38392__6417(.A (n_1683), .B (n_1147), .Y (n_1160));
  NOR2X1 g38388__5477(.A (n_1163), .B (n_770), .Y (n_1159));
  NOR2X1 g38391__2398(.A (n_1163), .B (n_834), .Y (n_1158));
  SDFFX1 DFF_237_Q_reg(.CK (CK), .D (n_1072), .SI (dft_sdi_13), .SE
       (SE), .Q (g1453), .QN (n_182));
  CLKINVX2 g38383(.A (n_1157), .Y (n_1486));
  SDFFX1 DFF_127_Q_reg(.CK (CK), .D (n_1093), .SI (g219), .SE (SE), .Q
       (g806), .QN (n_181));
  SDFFX1 DFF_296_Q_reg(.CK (CK), .D (n_1084), .SI (n_10), .SE (SE), .Q
       (g143), .QN (n_180));
  CLKINVX2 g38302(.A (n_1156), .Y (n_1211));
  OAI21X1 g38228__5107(.A0 (n_646), .A1 (n_1074), .B0 (g1834), .Y
       (n_1155));
  OAI21X1 g38126__6260(.A0 (n_845), .A1 (n_1076), .B0 (g611), .Y
       (n_1154));
  AND2X1 g38497__4319(.A (g109), .B (g1400), .Y (n_1153));
  CLKXOR2X1 g38259__8428(.A (g1828), .B (n_1073), .Y (n_1152));
  SDFFX1 DFF_269_Q_reg(.CK (CK), .D (n_1063), .SI (n_68), .SE (SE), .Q
       (g2648), .QN (n_179));
  AOI21X1 g38403__5526(.A0 (g1212), .A1 (n_1067), .B0 (n_1683), .Y
       (n_1157));
  SDFFX1 DFF_434_Q_reg(.CK (CK), .D (n_1071), .SI (n_1), .SE (SE), .Q
       (g4181), .QN (n_178));
  SDFFX1 DFF_279_Q_reg(.CK (CK), .D (n_1070), .SI (g1482), .SE (SE), .Q
       (g296), .QN (n_177));
  SDFFX1 DFF_215_Q_reg(.CK (CK), .D (g1356), .SI (n_211), .SE (SE), .Q
       (g1317), .QN (n_176));
  CLKINVX2 g38351(.A (n_1231), .Y (n_1151));
  OAI221X1 g38421__6783(.A0 (n_1146), .A1 (n_1149), .B0 (n_1083), .B1
       (n_1631), .C0 (n_1259), .Y (n_1150));
  NAND4X1 g38314__3680(.A (n_530), .B (n_1089), .C (n_1060), .D
       (n_1039), .Y (n_1148));
  NAND3X1 g38321__1617(.A (n_1097), .B (n_1096), .C (n_1212), .Y
       (n_1156));
  SDFFX1 DFF_347_Q_reg(.CK (CK), .D (n_1053), .SI (n_150), .SE (SE), .Q
       (g826), .QN (n_175));
  NAND2X1 g38374__2802(.A (g868), .B (g109), .Y (n_1566));
  SDFFX1 DFF_261_Q_reg(.CK (CK), .D (n_1055), .SI (n_248), .SE (SE), .Q
       (g617), .QN (n_174));
  XNOR2X1 g38465__1705(.A (n_1146), .B (g1462), .Y (n_1147));
  OR3X1 g38140__5122(.A (g704), .B (n_1085), .C (n_1138), .Y (n_1145));
  AOI21X1 g38092__8246(.A0 (n_1130), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1144));
  AOI21X1 g38093__7098(.A0 (n_1133), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1143));
  AOI21X1 g38094__6131(.A0 (n_1135), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1140));
  OR3X1 g38139__1881(.A (g686), .B (n_1103), .C (n_1138), .Y (n_1139));
  OR3X1 g38141__5115(.A (g668), .B (n_1109), .C (n_1138), .Y (n_1137));
  OR3X1 g38112__7482(.A (g731), .B (n_1135), .C (n_1138), .Y (n_1136));
  OR3X1 g38113__4733(.A (g677), .B (n_1133), .C (n_1138), .Y (n_1134));
  OR3X1 g38114__6161(.A (g713), .B (n_1105), .C (n_1138), .Y (n_1132));
  OR3X1 g38115__9315(.A (g695), .B (n_1130), .C (n_1138), .Y (n_1131));
  OR3X1 g38138__9945(.A (g722), .B (n_1107), .C (n_1138), .Y (n_1129));
  SDFFX1 DFF_389_Q_reg(.CK (CK), .D (n_1031), .SI (n_171), .SE (SE), .Q
       (g802), .QN (dft_sdo_21));
  SDFFX1 DFF_86_Q_reg(.CK (CK), .D (n_1013), .SI (n_146), .SE (SE), .Q
       (g736), .QN (n_172));
  SDFFX1 DFF_387_Q_reg(.CK (CK), .D (n_1020), .SI (n_131), .SE (SE), .Q
       (g818), .QN (n_171));
  SDFFX1 DFF_38_Q_reg(.CK (CK), .D (n_1030), .SI (g757), .SE (SE), .Q
       (g4180), .QN (n_170));
  SDFFX1 DFF_393_Q_reg(.CK (CK), .D (n_1018), .SI (n_91), .SE (SE), .Q
       (g810), .QN (n_169));
  SDFFX1 DFF_99_Q_reg(.CK (CK), .D (n_1036), .SI (g1470), .SE (SE), .Q
       (g822), .QN (n_168));
  OR2X2 g38484__2883(.A (g1212), .B (n_1683), .Y (n_1163));
  NOR2X1 g38150__2346(.A (n_1595), .B (n_1078), .Y (n_1128));
  NOR4X1 g38205__1666(.A (n_1239), .B (n_1068), .C (n_1293), .D
       (n_1052), .Y (n_1127));
  OR3X1 g38212__7410(.A (g658), .B (n_1079), .C (n_1138), .Y (n_1126));
  NOR2X1 g38281__6417(.A (n_1595), .B (n_1082), .Y (n_1125));
  OAI22X1 g38307__5477(.A0 (n_600), .A1 (n_1054), .B0 (n_701), .B1
       (n_1081), .Y (n_1124));
  NAND4X1 g38313__2398(.A (n_896), .B (n_965), .C (n_1065), .D
       (n_1001), .Y (n_1123));
  INVX1 g38349(.A (n_1102), .Y (n_1122));
  INVX1 g38348(.A (n_1101), .Y (n_1121));
  OAI211X1 g38422__5107(.A0 (n_1251), .A1 (n_1146), .B0 (n_503), .C0
       (n_1119), .Y (n_1120));
  SDFFX1 DFF_281_Q_reg(.CK (CK), .D (n_1016), .SI (n_119), .SE (SE), .Q
       (g700), .QN (n_167));
  SDFFX1 DFF_521_Q_reg(.CK (CK), .D (n_1010), .SI (n_75), .SE (SE), .Q
       (g691), .QN (n_166));
  SDFFX1 DFF_488_Q_reg(.CK (CK), .D (n_1021), .SI (g1380), .SE (SE), .Q
       (g673), .QN (n_165));
  SDFFX1 DFF_427_Q_reg(.CK (CK), .D (n_1017), .SI (n_345), .SE (SE), .Q
       (g727), .QN (n_164));
  SDFFX1 DFF_60_Q_reg(.CK (CK), .D (n_1014), .SI (n_115), .SE (SE), .Q
       (g682), .QN (n_163));
  SDFFX1 DFF_15_Q_reg(.CK (CK), .D (n_1009), .SI (n_374), .SE (SE), .Q
       (g709), .QN (n_162));
  SDFFX1 DFF_48_Q_reg(.CK (CK), .D (n_1015), .SI (n_264), .SE (SE), .Q
       (g718), .QN (n_161));
  SDFFX1 DFF_429_Q_reg(.CK (CK), .D (n_1026), .SI (n_50), .SE (SE), .Q
       (g798), .QN (n_160));
  SDFFX1 DFF_227_Q_reg(.CK (CK), .D (n_1033), .SI (n_142), .SE (SE), .Q
       (g794), .QN (n_159));
  CLKINVX2 g38353(.A (n_1118), .Y (n_1184));
  NAND4X1 g38377__6260(.A (n_1117), .B (n_700), .C (n_1116), .D
       (n_1115), .Y (n_1231));
  AOI21X1 g38164__4319(.A0 (n_1098), .A1 (n_985), .B0 (n_1113), .Y
       (n_1114));
  AOI21X1 g38125__8428(.A0 (n_1109), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1110));
  AOI21X1 g38124__5526(.A0 (n_1107), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1108));
  AOI21X1 g38091__6783(.A0 (n_1105), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1106));
  AOI21X1 g38122__3680(.A0 (n_1103), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1104));
  SDFFX1 DFF_182_Q_reg(.CK (CK), .D (n_998), .SI (dft_sdi_10), .SE
       (SE), .Q (g1400), .QN (n_158));
  SDFFX1 DFF_184_Q_reg(.CK (CK), .D (n_988), .SI (g309), .SE (SE), .Q
       (g814), .QN (n_157));
  NAND2X1 g38483__1617(.A (g869), .B (g109), .Y (n_1570));
  AOI222X1 g38356__2802(.A0 (g907), .A1 (n_1347), .B0 (n_1286), .B1
       (g296), .C0 (n_1265), .C1 (g272), .Y (n_1102));
  AOI222X1 g38355__1705(.A0 (g913), .A1 (n_1347), .B0 (n_1265), .B1
       (g278), .C0 (n_1222), .C1 (g38), .Y (n_1101));
  OAI211X1 g38223__5122(.A0 (n_628), .A1 (n_1075), .B0 (n_1099), .C0
       (n_1098), .Y (n_1100));
  SDFFX1 DFF_441_Q_reg(.CK (CK), .D (g874), .SI (n_361), .SE (SE), .Q
       (UNCONNECTED27), .QN (g868));
  AOI21X1 g38379__8246(.A0 (n_1097), .A1 (n_1096), .B0 (n_1115), .Y
       (n_1118));
  SDFFX1 DFF_528_Q_reg(.CK (CK), .D (n_977), .SI (n_237), .SE (SE), .Q
       (g1), .QN (n_156));
  SDFFX1 DFF_10_Q_reg(.CK (CK), .D (n_997), .SI (n_205), .SE (SE), .Q
       (g1558), .QN (n_155));
  SDFFX1 DFF_180_Q_reg(.CK (CK), .D (n_986), .SI (n_269), .SE (SE), .Q
       (g664), .QN (n_154));
  SDFFX1 DFF_223_Q_reg(.CK (CK), .D (n_987), .SI (n_220), .SE (SE), .Q
       (g1840), .QN (n_153));
  AOI22X1 g38431__7098(.A0 (n_1286), .A1 (g290), .B0 (n_1265), .B1
       (g266), .Y (n_1095));
  NOR2X1 g38180__6131(.A (n_1595), .B (n_1012), .Y (n_1094));
  CLKINVX1 g38461(.A (n_1061), .Y (n_1093));
  AOI22X1 g38473__1881(.A0 (n_1287), .A1 (g7), .B0 (n_1293), .B1
       (g1733), .Y (n_1092));
  NOR2X1 g38499__5115(.A (g631), .B (n_1209), .Y (n_1091));
  NOR2X1 g38500__7482(.A (g1849), .B (n_891), .Y (n_1090));
  AOI22X1 g38429__4733(.A0 (n_1286), .A1 (g299), .B0 (n_1265), .B1
       (g275), .Y (n_1089));
  AOI22X1 g38432__6161(.A0 (n_1265), .A1 (g284), .B0 (n_1087), .B1
       (g947), .Y (n_1088));
  AOI21X1 g38127__9315(.A0 (n_1085), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1086));
  NOR2X1 g38396__9945(.A (n_1683), .B (n_1040), .Y (n_1084));
  OAI21X1 g38556__2883(.A0 (g18), .A1 (n_1083), .B0 (n_1028), .Y
       (n_1111));
  SDFFX1 DFF_299_Q_reg(.CK (CK), .D (g1217), .SI (n_193), .SE (SE), .Q
       (g1212), .QN (n_152));
  SDFFX1 DFF_155_Q_reg(.CK (CK), .D (n_945), .SI (n_13), .SE (SE), .Q
       (g1950), .QN (n_151));
  NAND2X1 g38454__2346(.A (n_1204), .B (g9), .Y (n_1345));
  SDFFX1 DFF_346_Q_reg(.CK (CK), .D (n_956), .SI (n_81), .SE (SE), .Q
       (g1806), .QN (n_150));
  AOI22X1 g38357__1666(.A0 (g1828), .A1 (n_992), .B0 (g1822), .B1
       (n_1081), .Y (n_1082));
  AOI21X1 g38211__7410(.A0 (n_1079), .A1 (n_1142), .B0 (n_1141), .Y
       (n_1080));
  AOI22X1 g38217__6417(.A0 (g591), .A1 (n_972), .B0 (n_704), .B1
       (n_1011), .Y (n_1078));
  AOI22X1 g38433__5477(.A0 (n_1265), .A1 (g263), .B0 (g886), .B1
       (n_1050), .Y (n_1077));
  AOI211X1 g38206__2398(.A0 (n_971), .A1 (n_1075), .B0 (g617), .C0
       (n_1006), .Y (n_1076));
  AOI21X1 g38364__5107(.A0 (n_735), .A1 (n_1081), .B0 (g1840), .Y
       (n_1074));
  OAI21X1 g38365__6260(.A0 (n_618), .A1 (n_1081), .B0 (n_1116), .Y
       (n_1073));
  NOR2X1 g38389__4319(.A (n_1683), .B (n_1041), .Y (n_1072));
  SDFFX1 DFF_373_Q_reg(.CK (CK), .D (n_946), .SI (dft_sdi_21), .SE
       (SE), .Q (g1932), .QN (n_149));
  SDFFX1 DFF_339_Q_reg(.CK (CK), .D (n_948), .SI (dft_sdi_19), .SE
       (SE), .Q (g1923), .QN (n_148));
  SDFFX1 DFF_313_Q_reg(.CK (CK), .D (n_947), .SI (n_383), .SE (SE), .Q
       (g1941), .QN (n_147));
  SDFFX1 DFF_85_Q_reg(.CK (CK), .D (n_943), .SI (n_38), .SE (SE), .Q
       (g1896), .QN (n_146));
  SDFFX1 DFF_349_Q_reg(.CK (CK), .D (n_941), .SI (n_175), .SE (SE), .Q
       (g1887), .QN (n_145));
  SDFFX1 DFF_493_Q_reg(.CK (CK), .D (n_944), .SI (n_312), .SE (SE), .Q
       (g1905), .QN (n_144));
  SDFFX1 DFF_209_Q_reg(.CK (CK), .D (n_942), .SI (n_333), .SE (SE), .Q
       (g1914), .QN (n_143));
  CLKINVX2 g38385(.A (n_1115), .Y (n_1212));
  AOI211X1 g37998__8428(.A0 (n_951), .A1 (n_950), .B0 (n_1029), .C0
       (n_1062), .Y (n_1071));
  MX2X1 g38474__5526(.A (g139), .B (g296), .S0 (n_1602), .Y (n_1070));
  AOI222X1 g38475__6783(.A0 (n_1222), .A1 (g35), .B0 (n_1068), .B1
       (g1555), .C0 (n_1064), .C1 (g1531), .Y (n_1069));
  SDFFX1 DFF_226_Q_reg(.CK (CK), .D (n_1067), .SI (g318), .SE (SE), .Q
       (g1356), .QN (n_142));
  NAND2X1 g38498__3680(.A (n_1287), .B (g1), .Y (n_1066));
  AOI22X1 g38536__1617(.A0 (n_1239), .A1 (g1595), .B0 (n_1064), .B1
       (g1528), .Y (n_1065));
  CLKXOR2X1 g37991__2802(.A (n_1062), .B (g590), .Y (n_1063));
  OAI211X1 g38471__1705(.A0 (g806), .A1 (n_611), .B0 (n_1032), .C0
       (n_736), .Y (n_1061));
  AOI22X1 g38527__5122(.A0 (n_1171), .A1 (g1327), .B0 (n_1064), .B1
       (g1537), .Y (n_1060));
  AOI22X1 g38530__8246(.A0 (n_1296), .A1 (g1586), .B0 (n_1064), .B1
       (g1543), .Y (n_1059));
  AOI22X1 g38531__7098(.A0 (n_1068), .A1 (g1564), .B0 (n_1064), .B1
       (g1540), .Y (n_1058));
  AOI22X1 g38534__6131(.A0 (n_1068), .A1 (g1558), .B0 (n_1064), .B1
       (g1534), .Y (n_1057));
  AOI22X1 g38535__1881(.A0 (n_1064), .A1 (g1546), .B0 (g1191), .B1
       (n_1284), .Y (n_1056));
  SDFFX1 DFF_188_Q_reg(.CK (CK), .D (g875), .SI (n_238), .SE (SE), .Q
       (UNCONNECTED28), .QN (g869));
  SDFFX1 DFF_532_Q_reg(.CK (CK), .D (n_913), .SI (n_244), .SE (SE), .Q
       (g1878), .QN (dft_sdo_29));
  NOR2X1 g38182__5115(.A (n_1595), .B (n_981), .Y (n_1055));
  AOI21X1 g38387__7482(.A0 (g1822), .A1 (n_497), .B0 (n_1081), .Y
       (n_1054));
  NOR2X1 g38079__4733(.A (n_1035), .B (n_1002), .Y (n_1053));
  OR4X2 g38360__6161(.A (n_1051), .B (n_1050), .C (n_990), .D (n_963),
       .Y (n_1052));
  AOI222X1 g38420__9315(.A0 (n_1068), .A1 (g1549), .B0 (n_1293), .B1
       (g1721), .C0 (n_1064), .C1 (g1524), .Y (n_1049));
  OAI211X1 g38539__9945(.A0 (n_953), .A1 (n_952), .B0 (n_954), .C0
       (n_705), .Y (n_1048));
  XNOR2X1 g38572__2883(.A (g312), .B (g421), .Y (n_1047));
  AOI222X1 g38171__2346(.A0 (g722), .A1 (n_1024), .B0 (n_1046), .B1
       (n_1025), .C0 (g736), .C1 (n_1044), .Y (n_1135));
  AOI222X1 g38172__1666(.A0 (g686), .A1 (n_1023), .B0 (n_1045), .B1
       (n_1022), .C0 (g700), .C1 (n_1044), .Y (n_1130));
  AOI222X1 g38170__7410(.A0 (g668), .A1 (n_1008), .B0 (n_1043), .B1
       (n_1007), .C0 (g682), .C1 (n_1044), .Y (n_1133));
  SDFFX1 DFF_301_Q_reg(.CK (CK), .D (n_919), .SI (n_212), .SE (SE), .Q
       (g4179), .QN (n_140));
  AOI21X1 g38579__6417(.A0 (n_1595), .A1 (g1636), .B0 (n_1027), .Y
       (n_1146));
  NAND2X1 g38406__5477(.A (n_1116), .B (n_1081), .Y (n_1115));
  NAND4X1 g38278__2398(.A (n_1042), .B (n_610), .C (n_1099), .D
       (n_1004), .Y (n_1199));
  NAND2X1 g38245__5107(.A (n_1005), .B (n_1142), .Y (n_1138));
  CLKXOR2X1 g38464__6260(.A (g1453), .B (n_927), .Y (n_1041));
  CLKXOR2X1 g38467__4319(.A (g143), .B (n_931), .Y (n_1040));
  AOI222X1 g38477__8428(.A0 (n_1239), .A1 (g1604), .B0 (n_1068), .B1
       (g1561), .C0 (n_1296), .C1 (g1580), .Y (n_1039));
  AOI222X1 g38478__5526(.A0 (g892), .A1 (n_1050), .B0 (n_1037), .B1
       (g956), .C0 (n_1087), .C1 (g981), .Y (n_1038));
  NOR2X1 g38130__6783(.A (n_1035), .B (n_940), .Y (n_1036));
  INVX1 g38543(.A (n_1287), .Y (n_1034));
  SDFFX1 DFF_330_Q_reg(.CK (CK), .D (n_892), .SI (n_296), .SE (SE), .Q
       (UNCONNECTED29), .QN (g1849));
  SDFFX1 DFF_136_Q_reg(.CK (CK), .D (n_894), .SI (n_207), .SE (SE), .Q
       (UNCONNECTED30), .QN (g631));
  NAND2X1 g38588__3680(.A (n_1032), .B (g794), .Y (n_1033));
  AND2X1 g38591__1617(.A (n_564), .B (n_1032), .Y (n_1031));
  NOR2X1 g38035__2802(.A (n_1029), .B (n_964), .Y (n_1030));
  CLKINVX1 g38610(.A (n_1027), .Y (n_1028));
  OAI21X1 g38612__1705(.A0 (n_417), .A1 (n_563), .B0 (n_1032), .Y
       (n_1026));
  AOI211X1 g38220__5122(.A0 (g727), .A1 (n_1044), .B0 (n_1025), .C0
       (n_1024), .Y (n_1107));
  AOI211X1 g38184__8246(.A0 (g691), .A1 (n_1044), .B0 (n_1023), .C0
       (n_1022), .Y (n_1103));
  AOI222X1 g38169__7098(.A0 (g718), .A1 (n_1044), .B0 (n_689), .B1
       (n_967), .C0 (g704), .C1 (n_966), .Y (n_1105));
  NOR3X1 g38541__6131(.A (g42), .B (n_526), .C (n_991), .Y (n_1204));
  INVX1 g38252(.A (n_975), .Y (n_1021));
  AND2X1 g38231__1881(.A (n_865), .B (n_1032), .Y (n_1020));
  NOR2X1 g38234__5115(.A (g1909), .B (n_969), .Y (n_1019));
  AND2X1 g38283__7482(.A (n_743), .B (n_1032), .Y (n_1018));
  INVX1 g38247(.A (n_984), .Y (n_1017));
  INVX1 g38248(.A (n_979), .Y (n_1016));
  INVX1 g38249(.A (n_978), .Y (n_1015));
  INVX1 g38250(.A (n_989), .Y (n_1014));
  INVX1 g38251(.A (n_976), .Y (n_1013));
  AOI22X1 g38273__4733(.A0 (g605), .A1 (n_1011), .B0 (g599), .B1
       (n_1075), .Y (n_1012));
  INVX1 g38253(.A (n_974), .Y (n_1010));
  INVX1 g38254(.A (n_973), .Y (n_1009));
  AOI211X1 g38222__6161(.A0 (g673), .A1 (n_1044), .B0 (n_1008), .C0
       (n_1007), .Y (n_1109));
  INVX1 g38301(.A (n_1006), .Y (n_1098));
  SDFFX1 DFF_352_Q_reg(.CK (CK), .D (n_889), .SI (n_378), .SE (SE), .Q
       (g1845), .QN (n_139));
  SDFFX1 DFF_324_Q_reg(.CK (CK), .D (n_901), .SI (n_112), .SE (SE), .Q
       (g1796), .QN (dft_sdo_17));
  SDFFX1 DFF_104_Q_reg(.CK (CK), .D (n_898), .SI (n_60), .SE (SE), .Q
       (g1801), .QN (n_137));
  NOR2X1 g38246__9315(.A (n_1005), .B (n_1004), .Y (n_1141));
  AOI22X1 g38528__9945(.A0 (n_1296), .A1 (g1583), .B0 (n_1037), .B1
       (g965), .Y (n_1003));
  CLKXOR2X1 g38106__2883(.A (g826), .B (n_939), .Y (n_1002));
  AOI222X1 g38469__2346(.A0 (n_1037), .A1 (g953), .B0 (n_1087), .B1
       (g976), .C0 (g901), .C1 (n_1347), .Y (n_1001));
  AOI222X1 g38470__1666(.A0 (g919), .A1 (n_1347), .B0 (n_1222), .B1
       (g40), .C0 (n_1294), .C1 (g1311), .Y (n_1000));
  AOI222X1 g38476__7410(.A0 (n_1037), .A1 (g959), .B0 (n_1087), .B1
       (g986), .C0 (g895), .C1 (n_1050), .Y (n_999));
  NOR2X1 g38617__6417(.A (g248), .B (n_1683), .Y (n_998));
  OAI21X1 g38540__5477(.A0 (g1462), .A1 (n_1602), .B0 (n_639), .Y
       (n_997));
  AOI22X1 g38525__2398(.A0 (n_1239), .A1 (g1601), .B0 (g1179), .B1
       (n_1284), .Y (n_996));
  AOI22X1 g38526__5107(.A0 (n_1239), .A1 (g1598), .B0 (n_1296), .B1
       (g1574), .Y (n_995));
  SDFFX1 DFF_357_Q_reg(.CK (CK), .D (n_882), .SI (dft_sdi_20), .SE
       (SE), .Q (g874), .QN (n_136));
  AOI22X1 g38532__6260(.A0 (n_1037), .A1 (g968), .B0 (n_1087), .B1
       (g944), .Y (n_994));
  AOI22X1 g38533__4319(.A0 (n_1068), .A1 (g1552), .B0 (n_1296), .B1
       (g1571), .Y (n_993));
  SDFFX1 DFF_233_Q_reg(.CK (CK), .D (g1958), .SI (n_98), .SE (SE), .Q
       (UNCONNECTED31), .QN (g5816));
  NOR2X1 g38623__8428(.A (g248), .B (n_1595), .Y (n_1027));
  CLKINVX2 g38462(.A (n_992), .Y (n_1081));
  NOR2X1 g38561__5526(.A (n_876), .B (n_991), .Y (n_1287));
  AND2X2 g38511__6783(.A (n_888), .B (n_990), .Y (n_1286));
  AND2X2 g38514__3680(.A (g42), .B (n_990), .Y (n_1265));
  AOI22X1 g38264__1617(.A0 (g682), .A1 (n_983), .B0 (g673), .B1
       (n_982), .Y (n_989));
  NOR3X1 g38213__2802(.A (n_1035), .B (n_864), .C (n_728), .Y (n_988));
  NOR2X1 g38322__1705(.A (n_1595), .B (n_929), .Y (n_987));
  NAND3X1 g38225__5122(.A (n_1099), .B (n_870), .C (n_980), .Y (n_986));
  OAI21X1 g38235__8246(.A0 (n_968), .A1 (n_1075), .B0 (g622), .Y
       (n_985));
  AOI22X1 g38255__7098(.A0 (g727), .A1 (n_983), .B0 (g718), .B1
       (n_982), .Y (n_984));
  AOI22X1 g38261__6131(.A0 (n_804), .A1 (n_844), .B0 (g617), .B1
       (n_980), .Y (n_981));
  AOI22X1 g38262__1881(.A0 (g700), .A1 (n_983), .B0 (g691), .B1
       (n_982), .Y (n_979));
  AOI22X1 g38263__5115(.A0 (g718), .A1 (n_983), .B0 (g709), .B1
       (n_982), .Y (n_978));
  NOR2X1 g38168__7482(.A (n_1683), .B (n_914), .Y (n_977));
  AOI22X1 g38265__4733(.A0 (g736), .A1 (n_983), .B0 (g727), .B1
       (n_982), .Y (n_976));
  AOI22X1 g38267__6161(.A0 (g673), .A1 (n_983), .B0 (g664), .B1
       (n_982), .Y (n_975));
  AOI22X1 g38268__9315(.A0 (g691), .A1 (n_983), .B0 (g682), .B1
       (n_982), .Y (n_974));
  AOI22X1 g38269__9945(.A0 (g709), .A1 (n_983), .B0 (g700), .B1
       (n_982), .Y (n_973));
  OAI21X1 g38311__2883(.A0 (n_580), .A1 (n_971), .B0 (n_1011), .Y
       (n_972));
  INVX1 g38300(.A (n_969), .Y (n_970));
  NOR3X1 g38320__2346(.A (g622), .B (n_968), .C (n_1075), .Y (n_1006));
  AOI221X1 g38221__1666(.A0 (g709), .A1 (n_1044), .B0 (n_614), .B1
       (n_967), .C0 (n_966), .Y (n_1085));
  CLKINVX2 g38279(.A (n_1004), .Y (n_1142));
  AOI22X1 g38537__7410(.A0 (g889), .A1 (n_1050), .B0 (n_1222), .B1
       (g34), .Y (n_965));
  CLKXOR2X1 g38062__6417(.A (g4180), .B (n_842), .Y (n_964));
  NAND2X1 g38503__5477(.A (n_1309), .B (n_895), .Y (n_963));
  AOI22X1 g38520__2398(.A0 (n_1171), .A1 (g1321), .B0 (g1176), .B1
       (n_1284), .Y (n_962));
  AOI22X1 g38521__5107(.A0 (n_1171), .A1 (g1324), .B0 (n_1294), .B1
       (g1351), .Y (n_961));
  AOI22X1 g38522__6260(.A0 (g1194), .A1 (n_1320), .B0 (g1170), .B1
       (n_1284), .Y (n_960));
  AOI22X1 g38523__4319(.A0 (n_1294), .A1 (g1308), .B0 (n_1222), .B1
       (g39), .Y (n_959));
  AOI22X1 g38524__8428(.A0 (n_1171), .A1 (g1314), .B0 (n_1294), .B1
       (g1336), .Y (n_958));
  AOI22X1 g38529__5526(.A0 (n_1171), .A1 (g1318), .B0 (g1197), .B1
       (n_1320), .Y (n_957));
  OAI22X1 g38466__6783(.A0 (n_900), .A1 (n_857), .B0 (g1713), .B1
       (n_880), .Y (n_956));
  AOI22X1 g38538__3680(.A0 (g1182), .A1 (n_1284), .B0 (g910), .B1
       (n_1347), .Y (n_955));
  SDFFX1 DFF_137_Q_reg(.CK (CK), .D (n_860), .SI (g631), .SE (SE), .Q
       (g1217), .QN (n_135));
  NAND2X1 g38589__1617(.A (n_953), .B (n_952), .Y (n_954));
  SDFFX1 DFF_2_Q_reg(.CK (CK), .D (g255), .SI (n_213), .SE (SE), .Q
       (UNCONNECTED32), .QN (g312));
  NOR2X1 g38038__2802(.A (n_951), .B (n_950), .Y (n_1062));
  NOR2X1 g38485__1705(.A (n_1097), .B (n_899), .Y (n_992));
  SDFFX1 DFF_382_Q_reg(.CK (CK), .D (n_861), .SI (n_197), .SE (SE), .Q
       (g139), .QN (n_134));
  CLKINVX2 g38679(.A (n_1035), .Y (n_1032));
  INVX1 g38587(.A (n_949), .Y (n_1064));
  INVX1 g38408(.A (n_910), .Y (n_948));
  INVX1 g38407(.A (n_920), .Y (n_947));
  INVX1 g38410(.A (n_911), .Y (n_946));
  INVX1 g38413(.A (n_926), .Y (n_945));
  INVX1 g38412(.A (n_921), .Y (n_944));
  INVX1 g38411(.A (n_915), .Y (n_943));
  INVX1 g38414(.A (n_930), .Y (n_942));
  INVX1 g38409(.A (n_916), .Y (n_941));
  SDFFX1 DFF_196_Q_reg(.CK (CK), .D (n_843), .SI (n_274), .SE (SE), .Q
       (g654), .QN (n_133));
  OAI21X1 g38214__5122(.A0 (g822), .A1 (n_884), .B0 (n_939), .Y
       (n_940));
  SDFFX1 DFF_391_Q_reg(.CK (CK), .D (n_862), .SI (n_344), .SE (SE), .Q
       (g1524), .QN (n_132));
  AOI222X1 g38317__8246(.A0 (n_938), .A1 (n_934), .B0 (g1896), .B1
       (n_936), .C0 (g1882), .C1 (n_933), .Y (n_1182));
  AOI222X1 g38318__7098(.A0 (g1936), .A1 (n_907), .B0 (n_937), .B1
       (n_908), .C0 (g1950), .C1 (n_936), .Y (n_1180));
  AOI222X1 g38319__6131(.A0 (g1918), .A1 (n_905), .B0 (n_935), .B1
       (n_906), .C0 (g1932), .C1 (n_936), .Y (n_1185));
  AOI211X1 g38366__1881(.A0 (g1887), .A1 (n_936), .B0 (n_934), .C0
       (n_933), .Y (n_1188));
  SDFFX1 DFF_386_Q_reg(.CK (CK), .D (n_850), .SI (g1848), .SE (SE), .Q
       (g263), .QN (n_131));
  AOI222X1 g38316__5115(.A0 (g1914), .A1 (n_936), .B0 (n_932), .B1
       (n_902), .C0 (n_613), .C1 (n_903), .Y (n_969));
  NAND2X1 g38299__7482(.A (n_1099), .B (n_1075), .Y (n_1004));
  SDFFX1 DFF_247_Q_reg(.CK (CK), .D (n_849), .SI (n_185), .SE (SE), .Q
       (g4178), .QN (n_130));
  SDFFX1 DFF_72_Q_reg(.CK (CK), .D (n_846), .SI (n_339), .SE (SE), .Q
       (g639), .QN (n_129));
  CLKXOR2X1 g38577__4733(.A (g153), .B (n_848), .Y (n_931));
  AOI22X1 g38434__6161(.A0 (g1914), .A1 (n_925), .B0 (g1905), .B1
       (n_924), .Y (n_930));
  AOI22X1 g38435__9315(.A0 (n_928), .A1 (n_734), .B0 (g1840), .B1
       (n_912), .Y (n_929));
  SDFFX1 DFF_398_Q_reg(.CK (CK), .D (n_836), .SI (n_357), .SE (SE), .Q
       (g875), .QN (n_128));
  CLKXOR2X1 g38576__9945(.A (g1494), .B (n_851), .Y (n_927));
  AOI22X1 g38430__2883(.A0 (g1950), .A1 (n_925), .B0 (g1941), .B1
       (n_924), .Y (n_926));
  CLKXOR2X1 g38165__2346(.A (n_604), .B (n_922), .Y (n_923));
  AOI22X1 g38428__1666(.A0 (g1905), .A1 (n_925), .B0 (g1896), .B1
       (n_924), .Y (n_921));
  AOI22X1 g38423__7410(.A0 (g1941), .A1 (n_925), .B0 (g1932), .B1
       (n_924), .Y (n_920));
  SDFFX1 DFF_518_Q_reg(.CK (CK), .D (n_828), .SI (n_347), .SE (SE), .Q
       (g643), .QN (n_127));
  NOR2X1 g38085__6417(.A (n_1029), .B (n_867), .Y (n_919));
  NAND2X1 g38595__5477(.A (n_797), .B (n_917), .Y (n_991));
  OAI21X1 g38551__2398(.A0 (n_918), .A1 (g108), .B0 (g109), .Y
       (n_1067));
  SDFFX1 DFF_403_Q_reg(.CK (CK), .D (n_824), .SI (n_39), .SE (SE), .Q
       (g650), .QN (n_126));
  NAND2X1 g38609__5107(.A (n_874), .B (n_917), .Y (n_949));
  SDFFX1 DFF_76_Q_reg(.CK (CK), .D (n_840), .SI (dft_sdi_4), .SE (SE),
       .Q (UNCONNECTED33), .QN (g248));
  NOR3X1 g38578__6260(.A (g43), .B (n_525), .C (n_886), .Y (n_990));
  NAND3X1 g38719__4319(.A (g745), .B (g1957), .C (g109), .Y (n_1035));
  AOI22X1 g38425__8428(.A0 (g1887), .A1 (n_925), .B0 (g1878), .B1
       (n_924), .Y (n_916));
  AOI22X1 g38427__5526(.A0 (g1896), .A1 (n_925), .B0 (g1887), .B1
       (n_924), .Y (n_915));
  AOI21X1 g38177__6783(.A0 (n_1616), .A1 (n_847), .B0 (g1), .Y (n_914));
  NAND3X1 g38386__3680(.A (n_1116), .B (n_833), .C (n_912), .Y (n_913));
  AOI22X1 g38426__1617(.A0 (g1932), .A1 (n_925), .B0 (g1923), .B1
       (n_924), .Y (n_911));
  AOI22X1 g38424__2802(.A0 (g1923), .A1 (n_925), .B0 (g1914), .B1
       (n_924), .Y (n_910));
  MX2X1 g38218__1705(.A (n_852), .B (g1280), .S0 (g1284), .Y (n_909));
  AOI211X1 g38367__5122(.A0 (g1941), .A1 (n_936), .B0 (n_908), .C0
       (n_907), .Y (n_1175));
  AOI211X1 g38368__8246(.A0 (g1923), .A1 (n_936), .B0 (n_906), .C0
       (n_905), .Y (n_1173));
  SDFFX1 DFF_431_Q_reg(.CK (CK), .D (n_827), .SI (n_320), .SE (SE), .Q
       (g4172), .QN (n_125));
  AND2X1 g38291__7098(.A (n_967), .B (n_777), .Y (n_1025));
  SDFFX1 DFF_64_Q_reg(.CK (CK), .D (n_822), .SI (n_15), .SE (SE), .Q
       (g646), .QN (n_124));
  AND2X1 g38292__6131(.A (n_967), .B (n_904), .Y (n_1007));
  AND2X1 g38296__1881(.A (n_967), .B (n_547), .Y (n_1022));
  AOI221X1 g38370__5115(.A0 (g1905), .A1 (n_936), .B0 (n_546), .B1
       (n_903), .C0 (n_902), .Y (n_1178));
  CLKINVX2 g38352(.A (n_1075), .Y (n_1011));
  SDFFX1 DFF_30_Q_reg(.CK (CK), .D (n_825), .SI (n_355), .SE (SE), .Q
       (g4177), .QN (n_123));
  SDFFX1 DFF_143_Q_reg(.CK (CK), .D (n_831), .SI (g1365), .SE (SE), .Q
       (g1448), .QN (n_122));
  SDFFX1 DFF_174_Q_reg(.CK (CK), .D (n_821), .SI (n_44), .SE (SE), .Q
       (g1713), .QN (n_121));
  SDFFX1 DFF_111_Q_reg(.CK (CK), .D (n_818), .SI (n_359), .SE (SE), .Q
       (g1868), .QN (dft_sdo_5));
  OAI22X1 g38489__7482(.A0 (n_900), .A1 (n_837), .B0 (n_392), .B1
       (n_897), .Y (n_901));
  OAI221X1 g38490__4733(.A0 (n_937), .A1 (n_801), .B0 (g1936), .B1
       (n_810), .C0 (n_812), .Y (n_899));
  OAI22X1 g38515__6161(.A0 (n_788), .A1 (n_897), .B0 (n_900), .B1
       (n_795), .Y (n_898));
  NAND2X1 g38549__9315(.A (g925), .B (n_1051), .Y (n_896));
  NAND3X1 g38568__9945(.A (g45), .B (n_485), .C (n_879), .Y (n_895));
  NOR2X1 g38620__2883(.A (g630), .B (n_1209), .Y (n_894));
  INVX1 g38584(.A (n_1171), .Y (n_893));
  NOR2X1 g38619__2346(.A (g1848), .B (n_891), .Y (n_892));
  INVX1 g38586(.A (n_1284), .Y (n_890));
  NOR2X1 g38618__1666(.A (g1853), .B (n_891), .Y (n_889));
  SDFFX1 DFF_306_Q_reg(.CK (CK), .D (n_794), .SI (n_225), .SE (SE), .Q
       (UNCONNECTED34), .QN (g1462));
  NOR3X1 g38580__7410(.A (n_888), .B (n_887), .C (n_877), .Y (n_1293));
  INVX1 g38585(.A (n_1190), .Y (n_1037));
  NOR2X1 g38631__6417(.A (n_878), .B (n_886), .Y (n_1068));
  NOR2X1 g38604__5477(.A (n_875), .B (n_886), .Y (n_1239));
  NOR2X1 g38633__2398(.A (n_873), .B (n_886), .Y (n_1296));
  MX2X1 g38219__5107(.A (n_826), .B (g431), .S0 (g435), .Y (n_885));
  SDFFX1 DFF_280_Q_reg(.CK (CK), .D (n_803), .SI (n_177), .SE (SE), .Q
       (g1663), .QN (n_119));
  NAND2X1 g38086__6260(.A (g4180), .B (n_871), .Y (n_950));
  SDFFX1 DFF_18_Q_reg(.CK (CK), .D (n_816), .SI (n_90), .SE (SE), .Q
       (g1864), .QN (n_118));
  NAND2X1 g38709__4319(.A (g255), .B (g622), .Y (n_953));
  SDFFX1 DFF_159_Q_reg(.CK (CK), .D (n_807), .SI (g635), .SE (SE), .Q
       (g549), .QN (n_117));
  NAND2X1 g38237__8428(.A (g822), .B (n_884), .Y (n_939));
  NOR2X1 g38288__5526(.A (n_904), .B (n_883), .Y (n_1008));
  NOR2X1 g38294__6783(.A (n_648), .B (n_883), .Y (n_966));
  NOR2X1 g38295__3680(.A (n_544), .B (n_883), .Y (n_1023));
  NOR2X1 g38297__1617(.A (n_747), .B (n_883), .Y (n_1024));
  SDFFX1 DFF_141_Q_reg(.CK (CK), .D (n_815), .SI (n_88), .SE (SE), .Q
       (g1861), .QN (n_116));
  NAND2X1 g38329__2802(.A (g736), .B (n_982), .Y (n_980));
  SDFFX1 DFF_59_Q_reg(.CK (CK), .D (n_813), .SI (n_108), .SE (SE), .Q
       (g1786), .QN (n_115));
  SDFFX1 DFF_75_Q_reg(.CK (CK), .D (n_806), .SI (n_265), .SE (SE), .Q
       (g1791), .QN (dft_sdo_3));
  OAI211X1 g38378__1705(.A0 (n_866), .A1 (n_778), .B0 (n_791), .C0
       (n_835), .Y (n_1075));
  NOR2X1 g38376__5122(.A (n_1113), .B (n_982), .Y (n_983));
  OR4X2 g38493__8246(.A (g43), .B (g48), .C (g42), .D (n_798), .Y
       (n_882));
  SDFFX1 DFF_318_Q_reg(.CK (CK), .D (n_782), .SI (n_384), .SE (SE), .Q
       (g1958), .QN (n_113));
  CLKXOR2X1 g38463__7098(.A (g1027), .B (n_814), .Y (n_881));
  OAI21X1 g38565__6131(.A0 (n_631), .A1 (n_856), .B0 (g1806), .Y
       (n_880));
  AND2X1 g38450__1881(.A (n_903), .B (g1872), .Y (n_933));
  SDFFX1 DFF_322_Q_reg(.CK (CK), .D (n_780), .SI (n_230), .SE (SE), .Q
       (g1270), .QN (n_112));
  NOR2X1 g38704__5115(.A (n_859), .B (n_839), .Y (n_1317));
  CLKINVX1 g38677(.A (n_886), .Y (n_917));
  SDFFX1 DFF_355_Q_reg(.CK (CK), .D (n_764), .SI (n_216), .SE (SE), .Q
       (g1255), .QN (n_111));
  NAND2X1 g38606__7482(.A (n_598), .B (n_879), .Y (n_1190));
  SDFFX1 DFF_442_Q_reg(.CK (CK), .D (n_766), .SI (g868), .SE (SE), .Q
       (g1260), .QN (dft_sdo_24));
  NOR2X1 g38629__4733(.A (n_878), .B (n_877), .Y (n_1320));
  NOR3X1 g38628__6161(.A (n_876), .B (n_567), .C (n_853), .Y (n_1050));
  NOR2X1 g38605__9315(.A (n_875), .B (n_877), .Y (n_1171));
  AND2X2 g38607__9945(.A (n_874), .B (n_879), .Y (n_1347));
  NOR2X1 g38608__2883(.A (n_529), .B (n_877), .Y (n_1284));
  NOR2X1 g38632__2346(.A (n_873), .B (n_877), .Y (n_1294));
  NAND2X1 g38326__1666(.A (g664), .B (n_869), .Y (n_870));
  OAI21X1 g38323__7410(.A0 (g1227), .A1 (n_809), .B0 (n_690), .Y
       (n_868));
  OAI21X1 g38142__6417(.A0 (g4179), .A1 (n_819), .B0 (n_842), .Y
       (n_867));
  SDFFX1 DFF_89_Q_reg(.CK (CK), .D (g1957), .SI (g1362), .SE (SE), .Q
       (g745), .QN (n_109));
  SDFFX1 DFF_58_Q_reg(.CK (CK), .D (n_784), .SI (dft_sdi_3), .SE (SE),
       .Q (g1265), .QN (n_108));
  SDFFX1 DFF_510_Q_reg(.CK (CK), .D (n_760), .SI (n_51), .SE (SE), .Q
       (g1235), .QN (n_107));
  SDFFX1 DFF_32_Q_reg(.CK (CK), .D (n_753), .SI (n_123), .SE (SE), .Q
       (g1304), .QN (n_106));
  SDFFX1 DFF_498_Q_reg(.CK (CK), .D (n_762), .SI (n_57), .SE (SE), .Q
       (g1300), .QN (n_105));
  SDFFX1 DFF_250_Q_reg(.CK (CK), .D (n_767), .SI (n_283), .SE (SE), .Q
       (g1292), .QN (n_104));
  SDFFX1 DFF_202_Q_reg(.CK (CK), .D (n_759), .SI (n_61), .SE (SE), .Q
       (g1240), .QN (n_103));
  SDFFX1 DFF_334_Q_reg(.CK (CK), .D (n_771), .SI (n_209), .SE (SE), .Q
       (g1245), .QN (n_102));
  SDFFX1 DFF_486_Q_reg(.CK (CK), .D (n_761), .SI (n_80), .SE (SE), .Q
       (g1284), .QN (n_101));
  SDFFX1 DFF_401_Q_reg(.CK (CK), .D (n_769), .SI (n_370), .SE (SE), .Q
       (g1280), .QN (n_100));
  SDFFX1 DFF_61_Q_reg(.CK (CK), .D (n_768), .SI (n_163), .SE (SE), .Q
       (g1296), .QN (n_99));
  SDFFX1 DFF_231_Q_reg(.CK (CK), .D (n_756), .SI (n_326), .SE (SE), .Q
       (g1250), .QN (n_98));
  NOR2X1 g38375__5477(.A (n_866), .B (n_1044), .Y (n_967));
  ADDHX1 g38280__2398(.A (g818), .B (n_864), .CO (n_884), .S (n_865));
  NOR2X1 g38873__5107(.A (g750), .B (n_789), .Y (g4171));
  MX2X1 g38686__6260(.A (g1508), .B (g1524), .S0 (n_1602), .Y (n_862));
  SDFFX1 DFF_336_Q_reg(.CK (CK), .D (n_718), .SI (n_267), .SE (SE), .Q
       (UNCONNECTED35), .QN (g630));
  SDFFX1 DFF_489_Q_reg(.CK (CK), .D (n_746), .SI (n_165), .SE (SE), .Q
       (UNCONNECTED36), .QN (g1853));
  SDFFX1 DFF_385_Q_reg(.CK (CK), .D (n_737), .SI (n_240), .SE (SE), .Q
       (UNCONNECTED37), .QN (g1848));
  NOR2X1 g38621__4319(.A (n_1683), .B (n_802), .Y (n_861));
  OR3X1 g38614__8428(.A (g48), .B (n_859), .C (n_858), .Y (n_860));
  OR2X1 g38590__5526(.A (g1806), .B (n_856), .Y (n_857));
  NOR2X1 g38451__6783(.A (g1872), .B (n_854), .Y (n_934));
  NAND2X1 g38506__3680(.A (g1950), .B (n_924), .Y (n_912));
  NOR2X1 g38481__1617(.A (n_799), .B (n_855), .Y (n_907));
  NOR2X1 g38449__2802(.A (n_716), .B (n_855), .Y (n_905));
  NOR2X1 g38452__1705(.A (n_685), .B (n_854), .Y (n_906));
  NOR2X1 g38480__5122(.A (n_582), .B (n_854), .Y (n_902));
  NOR2X1 g38479__8246(.A (n_811), .B (n_854), .Y (n_908));
  SDFFX1 DFF_523_Q_reg(.CK (CK), .D (n_742), .SI (n_316), .SE (SE), .Q
       (g1776), .QN (n_97));
  NOR2X1 g38626__7098(.A (n_878), .B (n_853), .Y (n_1051));
  SDFFX1 DFF_332_Q_reg(.CK (CK), .D (n_741), .SI (n_317), .SE (SE), .Q
       (g1781), .QN (n_96));
  NOR2X1 g38630__6131(.A (n_873), .B (n_853), .Y (n_1087));
  NOR2X1 g38513__1881(.A (n_1414), .B (n_924), .Y (n_925));
  AOI21X1 g38285__5115(.A0 (dft_sdo_26), .A1 (n_750), .B0 (g1280), .Y
       (n_852));
  XNOR2X1 g38711__7482(.A (g1508), .B (g1499), .Y (n_851));
  OAI21X1 g38687__4733(.A0 (g182), .A1 (n_1602), .B0 (n_638), .Y
       (n_850));
  NOR2X1 g38151__6161(.A (n_1029), .B (n_790), .Y (n_849));
  CLKXOR2X1 g38710__9315(.A (g182), .B (g148), .Y (n_848));
  AND4X2 g38309__9945(.A (g1419), .B (g1515), .C (g1448), .D (n_785),
       .Y (n_847));
  OAI221X1 g38310__2883(.A0 (n_507), .A1 (n_845), .B0 (n_603), .B1
       (n_844), .C0 (n_1099), .Y (n_846));
  OAI21X1 g38362__2346(.A0 (n_683), .A1 (n_707), .B0 (n_793), .Y
       (n_843));
  SDFFX1 DFF_256_Q_reg(.CK (CK), .D (n_720), .SI (n_331), .SE (SE), .Q
       (g1561), .QN (n_95));
  SDFFX1 DFF_505_Q_reg(.CK (CK), .D (n_719), .SI (n_62), .SE (SE), .Q
       (g1528), .QN (n_94));
  CLKINVX2 g38163(.A (n_842), .Y (n_871));
  AOI21X1 g38277__1666(.A0 (n_396), .A1 (n_751), .B0 (n_457), .Y
       (n_922));
  AND2X1 g38701__7410(.A (g1361), .B (g3069), .Y (n_918));
  NAND2X1 g38702__6417(.A (g3007), .B (g876), .Y (n_1278));
  SDFFX1 DFF_270_Q_reg(.CK (CK), .D (n_726), .SI (n_179), .SE (SE), .Q
       (g255), .QN (dft_sdo_14));
  NOR2X1 g38330__5477(.A (g664), .B (n_841), .Y (n_1079));
  NAND2X1 g38369__2398(.A (n_792), .B (n_841), .Y (n_1005));
  SDFFX1 DFF_253_Q_reg(.CK (CK), .D (n_744), .SI (n_183), .SE (SE), .Q
       (g4176), .QN (n_92));
  NAND2X1 g38372__5107(.A (n_866), .B (n_841), .Y (n_883));
  NAND2X1 g38717__6260(.A (g48), .B (n_838), .Y (n_886));
  CLKINVX2 g38416(.A (n_869), .Y (n_982));
  NOR2X1 g38742__4319(.A (g1397), .B (n_1683), .Y (n_840));
  INVX1 g38725(.A (n_838), .Y (n_839));
  NAND3X1 g38613__8428(.A (g1791), .B (n_715), .C (n_830), .Y (n_837));
  NAND3X1 g38611__5526(.A (n_829), .B (n_528), .C (n_796), .Y (n_836));
  AOI22X1 g38519__6783(.A0 (g722), .A1 (n_748), .B0 (n_1046), .B1
       (n_866), .Y (n_835));
  CLKXOR2X1 g38518__3680(.A (g1223), .B (n_808), .Y (n_834));
  NAND2X1 g38496__1617(.A (g1878), .B (n_832), .Y (n_833));
  NOR2X1 g38495__2802(.A (n_1683), .B (n_781), .Y (n_831));
  SDFFX1 DFF_392_Q_reg(.CK (CK), .D (n_671), .SI (n_132), .SE (SE), .Q
       (g1577), .QN (n_91));
  SDFFX1 DFF_17_Q_reg(.CK (CK), .D (n_669), .SI (n_45), .SE (SE), .Q
       (g1574), .QN (n_90));
  SDFFX1 DFF_511_Q_reg(.CK (CK), .D (n_709), .SI (n_107), .SE (SE), .Q
       (g299), .QN (n_89));
  SDFFX1 DFF_140_Q_reg(.CK (CK), .D (n_714), .SI (g1466), .SE (SE), .Q
       (g1571), .QN (n_88));
  SDFFX1 DFF_254_Q_reg(.CK (CK), .D (n_712), .SI (n_92), .SE (SE), .Q
       (g1583), .QN (dft_sdo_13));
  SDFFX1 DFF_164_Q_reg(.CK (CK), .D (n_674), .SI (g1368), .SE (SE), .Q
       (g1531), .QN (n_86));
  SDFFX1 DFF_176_Q_reg(.CK (CK), .D (n_682), .SI (g333), .SE (SE), .Q
       (g269), .QN (n_85));
  SDFFX1 DFF_425_Q_reg(.CK (CK), .D (n_673), .SI (dft_sdi_24), .SE
       (SE), .Q (g1595), .QN (n_84));
  SDFFX1 DFF_42_Q_reg(.CK (CK), .D (n_672), .SI (n_354), .SE (SE), .Q
       (g1534), .QN (n_83));
  AOI21X1 g38624__1705(.A0 (n_820), .A1 (n_830), .B0 (n_686), .Y
       (n_897));
  NAND3X1 g38437__5122(.A (g617), .B (n_629), .C (n_844), .Y (n_869));
  CLKINVX1 g38678(.A (n_853), .Y (n_879));
  CLKINVX2 g38487(.A (n_855), .Y (n_903));
  SDFFX1 DFF_149_Q_reg(.CK (CK), .D (n_706), .SI (n_377), .SE (SE), .Q
       (g4175), .QN (n_82));
  OR2X2 g38716__8246(.A (n_829), .B (n_858), .Y (n_877));
  OR2X1 g38363__7098(.A (n_491), .B (n_823), .Y (n_828));
  AND2X1 g38868__6131(.A (n_492), .B (g1957), .Y (n_827));
  NOR2X1 g38286__1881(.A (g431), .B (n_749), .Y (n_826));
  NOR2X1 g38306__5115(.A (n_1029), .B (n_775), .Y (n_825));
  NOR2X1 g38325__7482(.A (n_708), .B (n_823), .Y (n_824));
  NOR2X1 g38361__4733(.A (n_596), .B (n_823), .Y (n_822));
  OAI22X1 g38801__6161(.A0 (g1710), .A1 (n_1149), .B0 (n_820), .B1
       (n_1631), .Y (n_821));
  SDFFX1 DFF_345_Q_reg(.CK (CK), .D (n_679), .SI (n_280), .SE (SE), .Q
       (g272), .QN (n_81));
  SDFFX1 DFF_485_Q_reg(.CK (CK), .D (n_711), .SI (n_30), .SE (SE), .Q
       (g266), .QN (n_80));
  SDFFX1 DFF_20_Q_reg(.CK (CK), .D (n_668), .SI (dft_sdi_1), .SE (SE),
       .Q (g1580), .QN (n_79));
  SDFFX1 DFF_456_Q_reg(.CK (CK), .D (n_697), .SI (n_206), .SE (SE), .Q
       (g1598), .QN (n_78));
  SDFFX1 DFF_218_Q_reg(.CK (CK), .D (n_670), .SI (dft_sdi_12), .SE
       (SE), .Q (g1601), .QN (n_77));
  SDFFX1 DFF_371_Q_reg(.CK (CK), .D (n_663), .SI (n_252), .SE (SE), .Q
       (g1592), .QN (n_76));
  SDFFX1 DFF_520_Q_reg(.CK (CK), .D (n_678), .SI (n_351), .SE (SE), .Q
       (g1567), .QN (n_75));
  SDFFX1 DFF_466_Q_reg(.CK (CK), .D (n_675), .SI (n_253), .SE (SE), .Q
       (g1586), .QN (n_74));
  SDFFX1 DFF_477_Q_reg(.CK (CK), .D (n_681), .SI (n_298), .SE (SE), .Q
       (g1607), .QN (n_73));
  NAND2X1 g38175__9315(.A (g4179), .B (n_819), .Y (n_842));
  SDFFX1 DFF_81_Q_reg(.CK (CK), .D (n_676), .SI (n_59), .SE (SE), .Q
       (g1604), .QN (n_72));
  SDFFX1 DFF_130_Q_reg(.CK (CK), .D (n_680), .SI (n_0), .SE (SE), .Q
       (g1564), .QN (n_71));
  SDFFX1 DFF_229_Q_reg(.CK (CK), .D (n_713), .SI (n_242), .SE (SE), .Q
       (g302), .QN (n_70));
  SDFFX1 DFF_138_Q_reg(.CK (CK), .D (n_677), .SI (n_135), .SE (SE), .Q
       (g1589), .QN (n_69));
  SDFFX1 DFF_268_Q_reg(.CK (CK), .D (n_696), .SI (n_11), .SE (SE), .Q
       (g1771), .QN (n_68));
  CLKINVX2 g38415(.A (n_841), .Y (n_1044));
  OAI21X1 g38492__9945(.A0 (n_616), .A1 (n_615), .B0 (n_817), .Y
       (n_818));
  AND2X1 g38501__2883(.A (n_817), .B (n_553), .Y (n_816));
  AND2X1 g38502__2346(.A (n_817), .B (n_449), .Y (n_815));
  CLKXOR2X1 g38575__1666(.A (g1023), .B (n_699), .Y (n_814));
  OAI22X1 g38574__7410(.A0 (n_900), .A1 (n_703), .B0 (n_385), .B1
       (n_805), .Y (n_813));
  OAI21X1 g38569__6417(.A0 (g1945), .A1 (n_811), .B0 (n_810), .Y
       (n_812));
  NOR2X1 g38548__5477(.A (n_386), .B (n_808), .Y (n_809));
  INVX1 g38675(.A (n_773), .Y (n_807));
  OAI22X1 g38566__2398(.A0 (n_692), .A1 (n_805), .B0 (n_900), .B1
       (n_693), .Y (n_806));
  NOR2X1 g38507__5107(.A (g1878), .B (n_1096), .Y (n_1169));
  NAND2X1 g38510__6260(.A (n_597), .B (n_1096), .Y (n_855));
  SDFFX1 DFF_112_Q_reg(.CK (CK), .D (n_630), .SI (dft_sdi_6), .SE (SE),
       .Q (g4173), .QN (n_67));
  NAND4X1 g38625__4319(.A (g47), .B (g48), .C (n_581), .D (n_665), .Y
       (n_1309));
  SDFFX1 DFF_372_Q_reg(.CK (CK), .D (n_632), .SI (n_76), .SE (SE), .Q
       (g1703), .QN (dft_sdo_20));
  OAI21X1 g38436__8428(.A0 (g617), .A1 (n_804), .B0 (n_844), .Y
       (n_841));
  NAND2X1 g38509__5526(.A (n_810), .B (n_1096), .Y (n_854));
  CLKINVX2 g38562(.A (n_832), .Y (n_924));
  INVX1 g38676(.A (n_787), .Y (n_803));
  CLKXOR2X1 g38683__6783(.A (n_725), .B (g166), .Y (n_802));
  NOR2X1 g38685__3680(.A (n_800), .B (n_799), .Y (n_801));
  NAND2X1 g38688__1617(.A (n_797), .B (n_796), .Y (n_798));
  OR2X1 g38693__2802(.A (g1801), .B (n_830), .Y (n_795));
  NOR2X1 g38695__1705(.A (n_1683), .B (n_733), .Y (n_794));
  INVX1 g38384(.A (n_823), .Y (n_793));
  INVX1 g38382(.A (n_791), .Y (n_792));
  SDFFX1 DFF_122_Q_reg(.CK (CK), .D (n_891), .SI (n_258), .SE (SE), .Q
       (g16), .QN (n_65));
  SDFFX1 DFF_262_Q_reg(.CK (CK), .D (n_1209), .SI (n_174), .SE (SE), .Q
       (g17), .QN (n_64));
  SDFFX1 DFF_93_Q_reg(.CK (CK), .D (g3007), .SI (n_268), .SE (SE), .Q
       (UNCONNECTED38), .QN (g876));
  SDFFX1 DFF_194_Q_reg(.CK (CK), .D (g3069), .SI (n_259), .SE (SE), .Q
       (UNCONNECTED39), .QN (g1361));
  CLKXOR2X1 g38276__5122(.A (g4178), .B (n_774), .Y (n_790));
  CLKINVX1 g38896(.A (g1957), .Y (n_789));
  NOR2X1 g38752__8246(.A (g47), .B (n_724), .Y (n_838));
  OR2X1 g38713__7098(.A (n_788), .B (n_830), .Y (n_856));
  NAND2X1 g38718__6131(.A (g48), .B (n_796), .Y (n_853));
  AOI222X1 g38697__1881(.A0 (n_772), .A1 (n_786), .B0 (g1663), .B1
       (n_1251), .C0 (g1718), .C1 (n_786), .Y (n_787));
  AND4X2 g38472__5115(.A (g1520), .B (g1440), .C (n_387), .D (n_656),
       .Y (n_785));
  OAI22X1 g38743__7482(.A0 (n_779), .A1 (n_783), .B0 (n_765), .B1
       (n_1384), .Y (n_784));
  AND4X2 g38571__4733(.A (g1806), .B (g1707), .C (g1690), .D (n_653),
       .Y (n_782));
  CLKXOR2X1 g38573__6161(.A (n_590), .B (n_654), .Y (n_781));
  OAI22X1 g38741__9315(.A0 (n_752), .A1 (n_783), .B0 (n_779), .B1
       (n_1384), .Y (n_780));
  AND2X1 g38593__9945(.A (n_777), .B (n_776), .Y (n_778));
  OAI21X1 g38419__2883(.A0 (g4177), .A1 (n_684), .B0 (n_774), .Y
       (n_775));
  AOI222X1 g38696__2346(.A0 (g1718), .A1 (n_1631), .B0 (n_772), .B1
       (n_1631), .C0 (g549), .C1 (n_1149), .Y (n_773));
  OAI22X1 g38738__1666(.A0 (n_754), .A1 (n_783), .B0 (n_758), .B1
       (n_1384), .Y (n_771));
  NOR2X1 g38698__7410(.A (g1231), .B (n_691), .Y (n_770));
  INVX1 g38721(.A (n_738), .Y (n_769));
  INVX1 g38722(.A (n_732), .Y (n_768));
  INVX1 g38723(.A (n_729), .Y (n_767));
  OAI22X1 g38726__6417(.A0 (n_765), .A1 (n_783), .B0 (n_763), .B1
       (n_1384), .Y (n_766));
  OAI22X1 g38730__5477(.A0 (n_763), .A1 (n_783), .B0 (n_755), .B1
       (n_1384), .Y (n_764));
  SDFFX1 DFF_407_Q_reg(.CK (CK), .D (n_620), .SI (n_311), .SE (SE), .Q
       (g4174), .QN (n_63));
  NAND3X1 g38581__2398(.A (g1840), .B (n_460), .C (n_928), .Y (n_832));
  CLKINVX2 g38563(.A (n_1096), .Y (n_936));
  INVX1 g38764(.A (n_722), .Y (n_762));
  INVX1 g38765(.A (n_721), .Y (n_761));
  OAI22X1 g38769__5107(.A0 (n_757), .A1 (n_783), .B0 (dft_sdo_26), .B1
       (n_1384), .Y (n_760));
  OAI22X1 g38770__6260(.A0 (n_758), .A1 (n_783), .B0 (n_757), .B1
       (n_1384), .Y (n_759));
  OAI22X1 g38771__4319(.A0 (n_755), .A1 (n_783), .B0 (n_754), .B1
       (n_1384), .Y (n_756));
  OAI22X1 g38785__8428(.A0 (n_398), .A1 (n_783), .B0 (n_752), .B1
       (n_1384), .Y (n_753));
  NOR4X1 g38354__5526(.A (g525), .B (g506), .C (g481), .D (n_661), .Y
       (n_751));
  NOR4X1 g38418__6783(.A (g1235), .B (g1260), .C (g1255), .D (n_659),
       .Y (n_750));
  NOR4X1 g38358__3680(.A (g386), .B (g411), .C (g406), .D (n_660), .Y
       (n_749));
  SDFFX1 DFF_504_Q_reg(.CK (CK), .D (n_607), .SI (n_251), .SE (SE), .Q
       (g1666), .QN (n_62));
  NOR2X1 g38315__1617(.A (n_390), .B (n_774), .Y (n_819));
  AOI21X1 g38400__2802(.A0 (n_501), .A1 (n_968), .B0 (n_845), .Y
       (n_791));
  SDFFX1 DFF_153_Q_reg(.CK (CK), .D (n_605), .SI (n_330), .SE (SE), .Q
       (UNCONNECTED40), .QN (g1397));
  SDFFX1 DFF_364_Q_reg(.CK (CK), .D (n_608), .SI (n_208), .SE (SE), .Q
       (UNCONNECTED41), .QN (g182));
  SDFFX1 DFF_201_Q_reg(.CK (CK), .D (n_606), .SI (n_250), .SE (SE), .Q
       (g1508), .QN (n_61));
  NAND2X1 g38758__1705(.A (g47), .B (n_723), .Y (n_858));
  NAND2X1 g38404__5122(.A (n_1099), .B (n_845), .Y (n_823));
  SDFFX1 DFF_103_Q_reg(.CK (CK), .D (n_627), .SI (g174), .SE (SE), .Q
       (g1766), .QN (n_60));
  SDFFX1 DFF_80_Q_reg(.CK (CK), .D (g756), .SI (n_348), .SE (SE), .Q
       (g1957), .QN (n_59));
  OR2X1 g38592__8246(.A (n_776), .B (n_747), .Y (n_748));
  INVX1 g38724(.A (n_745), .Y (n_746));
  NOR2X1 g38439__7098(.A (n_1029), .B (n_658), .Y (n_744));
  CLKXOR2X1 g38417__6131(.A (g810), .B (n_727), .Y (n_743));
  OAI22X1 g38700__1881(.A0 (n_557), .A1 (n_900), .B0 (n_465), .B1
       (n_740), .Y (n_742));
  OAI22X1 g38684__5115(.A0 (n_545), .A1 (n_740), .B0 (n_652), .B1
       (n_900), .Y (n_741));
  CLKXOR2X1 g38682__7482(.A (g1218), .B (n_694), .Y (n_739));
  AOI22X1 g38727__4733(.A0 (g1280), .A1 (n_731), .B0 (g1284), .B1
       (n_730), .Y (n_738));
  OR2X1 g38733__6161(.A (g1845), .B (n_891), .Y (n_737));
  OR3X1 g38751__9315(.A (g31), .B (g30), .C (n_662), .Y (g9451));
  SDFFX1 DFF_234_Q_reg(.CK (CK), .D (n_593), .SI (g5816), .SE (SE), .Q
       (g1032), .QN (n_58));
  NOR2X1 g38457__9945(.A (n_594), .B (n_736), .Y (n_864));
  SDFFX1 DFF_497_Q_reg(.CK (CK), .D (n_576), .SI (n_263), .SE (SE), .Q
       (g991), .QN (n_57));
  OAI21X1 g38554__2883(.A0 (n_502), .A1 (n_735), .B0 (n_928), .Y
       (n_1097));
  SDFFX1 DFF_115_Q_reg(.CK (CK), .D (n_574), .SI (n_289), .SE (SE), .Q
       (g1015), .QN (n_56));
  SDFFX1 DFF_414_Q_reg(.CK (CK), .D (n_572), .SI (n_53), .SE (SE), .Q
       (g1003), .QN (n_55));
  SDFFX1 DFF_108_Q_reg(.CK (CK), .D (n_577), .SI (n_380), .SE (SE), .Q
       (g1007), .QN (n_54));
  SDFFX1 DFF_413_Q_reg(.CK (CK), .D (n_570), .SI (n_7), .SE (SE), .Q
       (g1027), .QN (n_53));
  NOR2X1 g38559__2346(.A (n_1414), .B (n_928), .Y (n_817));
  CLKINVX2 g38438(.A (n_845), .Y (n_844));
  OAI21X1 g38582__1666(.A0 (g1840), .A1 (n_734), .B0 (n_928), .Y
       (n_1096));
  SDFFX1 DFF_113_Q_reg(.CK (CK), .D (n_575), .SI (n_67), .SE (SE), .Q
       (g1718), .QN (n_52));
  CLKXOR2X1 g38800__7410(.A (dft_sdo_8), .B (n_772), .Y (n_733));
  AOI22X1 g38737__6417(.A0 (g1296), .A1 (n_731), .B0 (g1300), .B1
       (n_730), .Y (n_732));
  AOI22X1 g38749__5477(.A0 (g1292), .A1 (n_731), .B0 (g1296), .B1
       (n_730), .Y (n_729));
  AOI21X1 g38305__2398(.A0 (g810), .A1 (n_727), .B0 (g814), .Y (n_728));
  SDFFX1 DFF_471_Q_reg(.CK (CK), .D (n_633), .SI (n_286), .SE (SE), .Q
       (UNCONNECTED42), .QN (g1710));
  INVX1 g38849(.A (n_725), .Y (n_726));
  INVX1 g38805(.A (n_723), .Y (n_724));
  AOI22X1 g38767__5107(.A0 (g1300), .A1 (n_731), .B0 (g1304), .B1
       (n_730), .Y (n_722));
  AOI22X1 g38768__6260(.A0 (g1284), .A1 (n_731), .B0 (g1292), .B1
       (n_730), .Y (n_721));
  OAI21X1 g38772__4319(.A0 (dft_sdo_8), .A1 (n_1602), .B0 (n_636), .Y
       (n_720));
  OAI21X1 g38777__8428(.A0 (g1504), .A1 (n_1602), .B0 (n_635), .Y
       (n_719));
  OR2X1 g38734__5526(.A (g627), .B (n_1209), .Y (n_718));
  SDFFX1 DFF_509_Q_reg(.CK (CK), .D (n_591), .SI (g127), .SE (SE), .Q
       (g1618), .QN (n_51));
  OR3X1 g38755__6783(.A (n_935), .B (n_717), .C (n_716), .Y (n_799));
  NAND2X1 g38759__3680(.A (g1218), .B (n_657), .Y (n_808));
  SDFFX1 DFF_428_Q_reg(.CK (CK), .D (n_569), .SI (n_164), .SE (SE), .Q
       (g999), .QN (n_50));
  NOR2X1 g38757__1617(.A (g47), .B (n_664), .Y (n_796));
  SDFFX1 DFF_192_Q_reg(.CK (CK), .D (n_578), .SI (n_219), .SE (SE), .Q
       (g1023), .QN (n_49));
  SDFFX1 DFF_87_Q_reg(.CK (CK), .D (n_568), .SI (n_172), .SE (SE), .Q
       (g1019), .QN (n_48));
  NAND3X1 g38762__2802(.A (g1796), .B (g1791), .C (n_715), .Y (n_830));
  SDFFX1 DFF_167_Q_reg(.CK (CK), .D (n_573), .SI (n_226), .SE (SE), .Q
       (UNCONNECTED43), .QN (g1011));
  SDFFX1 DFF_515_Q_reg(.CK (CK), .D (n_571), .SI (n_218), .SE (SE), .Q
       (g995), .QN (n_47));
  MX2X1 g38780__1705(.A (g1520), .B (g1571), .S0 (n_1602), .Y (n_714));
  MX2X1 g38779__5122(.A (g143), .B (g302), .S0 (n_1602), .Y (n_713));
  MX2X1 g38778__8246(.A (g1424), .B (g1583), .S0 (n_1602), .Y (n_712));
  MX2X1 g38776__7098(.A (g178), .B (g266), .S0 (n_1602), .Y (n_711));
  CLKXOR2X1 g38775__6131(.A (g516), .B (n_584), .Y (n_710));
  MX2X1 g38774__1881(.A (g166), .B (g299), .S0 (n_1602), .Y (n_709));
  AOI21X1 g38564__5115(.A0 (g650), .A1 (n_612), .B0 (n_707), .Y
       (n_708));
  NOR2X1 g38616__7482(.A (n_1029), .B (n_625), .Y (n_706));
  OR4X1 g38689__4733(.A (n_704), .B (n_602), .C (n_609), .D (n_804), .Y
       (n_705));
  NAND3X1 g38690__6161(.A (g1781), .B (n_566), .C (n_687), .Y (n_703));
  NAND4X1 g38691__9315(.A (n_701), .B (n_601), .C (n_700), .D (n_592),
       .Y (n_702));
  CLKXOR2X1 g38703__9945(.A (n_552), .B (n_589), .Y (n_699));
  CLKXOR2X1 g38773__2883(.A (g501), .B (n_586), .Y (n_698));
  MX2X1 g38766__2346(.A (g1436), .B (g1598), .S0 (n_1602), .Y (n_697));
  OAI21X1 g38740__1666(.A0 (n_440), .A1 (n_900), .B0 (n_619), .Y
       (n_696));
  NAND2X1 g38735__7410(.A (g1227), .B (n_694), .Y (n_695));
  NAND2X1 g38736__6417(.A (n_692), .B (n_715), .Y (n_693));
  NOR2X1 g38739__5477(.A (n_690), .B (n_694), .Y (n_691));
  NAND2X1 g38750__2398(.A (g1850), .B (n_647), .Y (n_745));
  CLKAND2X2 g38712__5107(.A (n_689), .B (n_688), .Y (n_777));
  AOI21X1 g38708__6260(.A0 (n_820), .A1 (n_687), .B0 (n_686), .Y
       (n_805));
  OR3X1 g38705__4319(.A (g1918), .B (g1927), .C (n_685), .Y (n_811));
  SDFFX1 DFF_292_Q_reg(.CK (CK), .D (n_534), .SI (dft_sdi_16), .SE
       (SE), .Q (g1071), .QN (n_46));
  SDFFX1 DFF_16_Q_reg(.CK (CK), .D (n_527), .SI (n_162), .SE (SE), .Q
       (g1092), .QN (n_45));
  SDFFX1 DFF_173_Q_reg(.CK (CK), .D (n_539), .SI (n_241), .SE (SE), .Q
       (g1080), .QN (n_44));
  SDFFX1 DFF_290_Q_reg(.CK (CK), .D (n_559), .SI (n_371), .SE (SE), .Q
       (g1089), .QN (dft_sdo_15));
  NAND2X1 g38482__8428(.A (g4177), .B (n_684), .Y (n_774));
  NAND2X1 g38460__5526(.A (n_683), .B (n_707), .Y (n_845));
  MX2X1 g38792__6783(.A (g148), .B (g269), .S0 (n_1602), .Y (n_682));
  MX2X1 g38783__3680(.A (g1448), .B (g1607), .S0 (n_1602), .Y (n_681));
  MX2X1 g38784__1617(.A (g1453), .B (g1564), .S0 (n_1602), .Y (n_680));
  MX2X1 g38786__2802(.A (g153), .B (g272), .S0 (n_1602), .Y (n_679));
  MX2X1 g38787__1705(.A (g1415), .B (g1567), .S0 (n_1602), .Y (n_678));
  MX2X1 g38788__5122(.A (g1428), .B (g1589), .S0 (n_1602), .Y (n_677));
  MX2X1 g38789__8246(.A (g1444), .B (g1604), .S0 (n_1602), .Y (n_676));
  MX2X1 g38790__7098(.A (g1407), .B (g1586), .S0 (n_1602), .Y (n_675));
  MX2X1 g38791__6131(.A (g1499), .B (g1531), .S0 (n_1602), .Y (n_674));
  MX2X1 g38782__1881(.A (g1432), .B (g1595), .S0 (n_1602), .Y (n_673));
  MX2X1 g38793__5115(.A (g1494), .B (g1534), .S0 (n_1602), .Y (n_672));
  MX2X1 g38794__7482(.A (g1419), .B (g1577), .S0 (n_1602), .Y (n_671));
  MX2X1 g38795__4733(.A (g1440), .B (g1601), .S0 (n_1602), .Y (n_670));
  MX2X1 g38796__6161(.A (g1515), .B (g1574), .S0 (n_1602), .Y (n_669));
  MX2X1 g38797__9315(.A (g1411), .B (g1580), .S0 (n_1602), .Y (n_668));
  CLKXOR2X1 g38799__9945(.A (g476), .B (n_587), .Y (n_667));
  CLKXOR2X1 g38802__2883(.A (g491), .B (n_588), .Y (n_666));
  CLKINVX1 g38847(.A (n_664), .Y (n_665));
  MX2X1 g38781__2346(.A (g1403), .B (g1592), .S0 (n_1602), .Y (n_663));
  SDFFX1 DFF_170_Q_reg(.CK (CK), .D (n_531), .SI (n_27), .SE (SE), .Q
       (g1074), .QN (n_42));
  SDFFX1 DFF_94_Q_reg(.CK (CK), .D (n_540), .SI (g876), .SE (SE), .Q
       (g1086), .QN (dft_sdo_4));
  AOI21X1 g38886__1666(.A0 (n_1595), .A1 (g549), .B0 (n_772), .Y
       (n_725));
  SDFFX1 DFF_56_Q_reg(.CK (CK), .D (n_533), .SI (n_9), .SE (SE), .Q
       (g1095), .QN (n_40));
  SDFFX1 DFF_402_Q_reg(.CK (CK), .D (n_532), .SI (n_100), .SE (SE), .Q
       (g1083), .QN (n_39));
  SDFFX1 DFF_82_Q_reg(.CK (CK), .D (n_535), .SI (n_72), .SE (SE), .Q
       (g1098), .QN (n_38));
  SDFFX1 DFF_27_Q_reg(.CK (CK), .D (n_536), .SI (n_360), .SE (SE), .Q
       (g1077), .QN (n_37));
  SDFFX1 DFF_376_Q_reg(.CK (CK), .D (n_561), .SI (n_337), .SE (SE), .Q
       (g1068), .QN (n_36));
  NOR2X1 g38812__7410(.A (g46), .B (n_662), .Y (n_723));
  OR4X1 g38516__6417(.A (g476), .B (g491), .C (g516), .D (n_555), .Y
       (n_661));
  OR4X1 g38517__5477(.A (g421), .B (g416), .C (g391), .D (n_556), .Y
       (n_660));
  OR4X1 g38567__2398(.A (g1245), .B (g1250), .C (g1270), .D (n_554), .Y
       (n_659));
  CLKXOR2X1 g38570__5107(.A (g4176), .B (n_624), .Y (n_658));
  CLKINVX2 g38850(.A (n_694), .Y (n_657));
  AND4X2 g38615__6260(.A (g1428), .B (g1432), .C (n_432), .D (n_550),
       .Y (n_656));
  NAND2X1 g38807__4319(.A (g1537), .B (n_1602), .Y (n_655));
  CLKXOR2X1 g38706__8428(.A (g1448), .B (n_551), .Y (n_654));
  NOR3X1 g38745__5526(.A (n_518), .B (n_517), .C (n_652), .Y (n_653));
  CLKXOR2X1 g38803__6783(.A (n_650), .B (n_560), .Y (n_651));
  CLKINVX2 g38486(.A (n_727), .Y (n_736));
  OR3X1 g38707__3680(.A (n_688), .B (n_649), .C (n_648), .Y (n_747));
  SDFFX1 DFF_53_Q_reg(.CK (CK), .D (n_522), .SI (n_375), .SE (SE), .Q
       (g3007), .QN (n_35));
  SDFFX1 DFF_328_Q_reg(.CK (CK), .D (n_521), .SI (n_276), .SE (SE), .Q
       (g3069), .QN (n_34));
  CLKINVX2 g38852(.A (n_647), .Y (n_891));
  SDFFX1 DFF_276_Q_reg(.CK (CK), .D (n_516), .SI (g1959), .SE (SE), .Q
       (g1690), .QN (n_33));
  CLKINVX2 g38583(.A (n_646), .Y (n_928));
  NAND2X1 g38866__1617(.A (g293), .B (n_1602), .Y (n_645));
  NAND2X1 g38856__2802(.A (g281), .B (n_1602), .Y (n_644));
  NAND2X1 g38858__1705(.A (g1543), .B (n_1602), .Y (n_643));
  NAND2X1 g38859__5122(.A (g278), .B (n_1602), .Y (n_642));
  NAND2X1 g38860__8246(.A (g287), .B (n_1602), .Y (n_641));
  NAND2X1 g38861__7098(.A (g1552), .B (n_1602), .Y (n_640));
  NAND2X1 g38863__6131(.A (g1558), .B (n_1602), .Y (n_639));
  NAND2X1 g38864__1881(.A (g263), .B (n_1602), .Y (n_638));
  NAND2X1 g38865__5115(.A (g1555), .B (n_1602), .Y (n_637));
  NAND2X1 g38855__7482(.A (g1561), .B (n_1602), .Y (n_636));
  NAND2X1 g38867__4733(.A (g1528), .B (n_1602), .Y (n_635));
  NOR2X1 g38913__6161(.A (g1696), .B (n_633), .Y (g6842));
  AOI21X1 g38943__9315(.A0 (n_631), .A1 (n_1251), .B0 (n_633), .Y
       (n_632));
  NOR2X1 g38908__9945(.A (n_1029), .B (g4173), .Y (n_630));
  NAND2X1 g38883__2883(.A (g46), .B (n_599), .Y (n_664));
  SDFFX1 DFF_380_Q_reg(.CK (CK), .D (n_520), .SI (n_291), .SE (SE), .Q
       (g9), .QN (n_32));
  OAI21X1 g38892__2346(.A0 (g591), .A1 (n_629), .B0 (n_1099), .Y
       (n_1209));
  CLKINVX2 g38897(.A (n_731), .Y (n_783));
  AOI211X1 g38874__1666(.A0 (g599), .A1 (n_499), .B0 (n_488), .C0
       (n_579), .Y (n_628));
  OAI221X1 g38872__7410(.A0 (g1766), .A1 (n_631), .B0 (n_439), .B1
       (n_626), .C0 (n_820), .Y (n_627));
  OAI21X1 g38747__6417(.A0 (g4175), .A1 (n_543), .B0 (n_624), .Y
       (n_625));
  CLKXOR2X1 g38862__5477(.A (g496), .B (n_495), .Y (n_623));
  CLKXOR2X1 g38798__2398(.A (g511), .B (n_512), .Y (n_622));
  XNOR2X1 g38804__5107(.A (g486), .B (n_514), .Y (n_621));
  AND2X1 g38808__6260(.A (n_483), .B (n_565), .Y (n_620));
  OAI21X1 g38857__4319(.A0 (n_420), .A1 (n_686), .B0 (g1771), .Y
       (n_619));
  AOI211X1 g38853__8428(.A0 (g1822), .A1 (n_486), .B0 (n_489), .C0
       (n_583), .Y (n_618));
  CLKXOR2X1 g38854__5526(.A (g506), .B (n_493), .Y (n_617));
  NAND2X1 g38603__6783(.A (n_616), .B (n_615), .Y (n_646));
  AND2X1 g38753__3680(.A (n_614), .B (n_649), .Y (n_689));
  NAND2X1 g38811__1617(.A (g1909), .B (n_613), .Y (n_716));
  NOR2X1 g38622__2802(.A (n_402), .B (n_624), .Y (n_684));
  NOR2X1 g38599__1705(.A (g650), .B (n_612), .Y (n_707));
  CLKAND2X2 g38627__5122(.A (g806), .B (n_611), .Y (n_727));
  CLKINVX2 g38851(.A (n_687), .Y (n_715));
  INVX1 g38933(.A (n_609), .Y (n_610));
  AND2X1 g38900__8246(.A (g109), .B (g178), .Y (n_608));
  OAI21X1 g38907__7098(.A0 (n_471), .A1 (n_786), .B0 (n_1119), .Y
       (n_607));
  NOR2X1 g38909__6131(.A (g1504), .B (n_1683), .Y (n_606));
  NOR2X1 g38914__1881(.A (g192), .B (n_1683), .Y (n_605));
  NOR2X1 g38918__5115(.A (g471), .B (n_542), .Y (n_604));
  SDFFX1 DFF_68_Q_reg(.CK (CK), .D (g755), .SI (g1371), .SE (SE), .Q
       (g756), .QN (n_31));
  AOI21X1 g38877__7482(.A0 (n_820), .A1 (n_508), .B0 (n_686), .Y
       (n_740));
  AOI22X1 g38884__4733(.A0 (n_603), .A1 (n_602), .B0 (g639), .B1
       (n_704), .Y (n_952));
  OAI22X1 g38875__6161(.A0 (g1857), .A1 (n_601), .B0 (n_505), .B1
       (n_701), .Y (n_1281));
  AOI21X1 g38891__9315(.A0 (g1834), .A1 (n_600), .B0 (n_1414), .Y
       (n_647));
  CLKINVX1 g38894(.A (n_599), .Y (n_662));
  INVX1 g38934(.A (n_598), .Y (n_875));
  CLKINVX2 g38895(.A (n_597), .Y (n_810));
  NAND2X1 g38889__9945(.A (n_730), .B (n_1360), .Y (n_694));
  NOR2X1 g38929__2883(.A (g192), .B (n_1595), .Y (n_772));
  NOR2X1 g38931__2346(.A (n_1683), .B (n_730), .Y (n_731));
  AOI21X1 g38746__1666(.A0 (g646), .A1 (n_498), .B0 (n_549), .Y
       (n_596));
  AOI211X1 g38699__7410(.A0 (n_424), .A1 (n_594), .B0 (n_400), .C0
       (n_476), .Y (n_595));
  MX2X1 g38955__6417(.A (g1077), .B (g1032), .S0 (n_1149), .Y (n_593));
  INVX1 g38848(.A (n_734), .Y (n_592));
  MX2X1 g38869__5477(.A (n_590), .B (g1618), .S0 (n_1149), .Y (n_591));
  CLKXOR2X1 g38880__2398(.A (n_450), .B (n_482), .Y (n_589));
  NAND2X1 g38923__5107(.A (n_511), .B (n_585), .Y (n_588));
  NAND2X1 g38919__6260(.A (g471), .B (n_510), .Y (n_587));
  NAND2X1 g38921__4319(.A (g461), .B (n_585), .Y (n_586));
  NAND2X1 g38922__8428(.A (g471), .B (n_541), .Y (n_584));
  SDFFX1 DFF_484_Q_reg(.CK (CK), .D (n_438), .SI (n_329), .SE (SE), .Q
       (g1374), .QN (n_30));
  OR2X2 g38928__5526(.A (n_468), .B (n_583), .Y (n_597));
  OR3X1 g38881__6783(.A (g1900), .B (g1909), .C (n_582), .Y (n_685));
  AOI21X1 g38924__3680(.A0 (n_412), .A1 (n_1222), .B0 (g41), .Y
       (n_599));
  SDFFX1 DFF_77_Q_reg(.CK (CK), .D (n_437), .SI (g248), .SE (SE), .Q
       (g1707), .QN (n_29));
  INVX1 g38935(.A (n_581), .Y (n_878));
  OR2X1 g38927__1617(.A (n_580), .B (n_579), .Y (n_866));
  CLKINVX2 g38937(.A (n_1113), .Y (n_1099));
  INVX4 g38898(.A (n_562), .Y (n_1602));
  MX2X1 g38953__2802(.A (g1071), .B (g1023), .S0 (n_1149), .Y (n_578));
  MX2X1 g38938__1705(.A (g1095), .B (g1007), .S0 (n_1149), .Y (n_577));
  MX2X1 g38945__5122(.A (g1083), .B (g991), .S0 (n_1149), .Y (n_576));
  OAI22X1 g38946__8246(.A0 (n_820), .A1 (n_1149), .B0 (n_484), .B1
       (n_1631), .Y (n_575));
  MX2X1 g38949__7098(.A (g1074), .B (g1015), .S0 (n_1149), .Y (n_574));
  OAI22X1 g38947__6131(.A0 (n_389), .A1 (n_1149), .B0 (g1011), .B1
       (n_1631), .Y (n_573));
  MX2X1 g38948__1881(.A (g1086), .B (g1003), .S0 (n_1149), .Y (n_572));
  MX2X1 g38950__5115(.A (g1080), .B (g995), .S0 (n_1149), .Y (n_571));
  MX2X1 g38952__7482(.A (g1068), .B (g1027), .S0 (n_1149), .Y (n_570));
  MX2X1 g38956__4733(.A (g1089), .B (g999), .S0 (n_1149), .Y (n_569));
  MX2X1 g38954__6161(.A (g1098), .B (g1019), .S0 (n_1149), .Y (n_568));
  OAI21X1 g38964__9315(.A0 (g605), .A1 (n_580), .B0 (n_968), .Y
       (n_609));
  NOR3X1 g38968__9945(.A (g43), .B (g42), .C (n_567), .Y (n_598));
  SDFFX1 DFF_165_Q_reg(.CK (CK), .D (n_435), .SI (n_86), .SE (SE), .Q
       (UNCONNECTED44), .QN (dft_sdo_8));
  NAND3X1 g38890__2883(.A (g1781), .B (g1786), .C (n_566), .Y (n_687));
  NAND2X1 g39003__2346(.A (g1700), .B (g1959), .Y (n_633));
  SDFFX1 DFF_90_Q_reg(.CK (CK), .D (n_433), .SI (n_109), .SE (SE), .Q
       (g1419), .QN (n_28));
  CLKINVX2 g38936(.A (n_1414), .Y (n_1116));
  CLKINVX2 g39028(.A (n_565), .Y (n_1029));
  ADDHX1 g38634__1666(.A (g802), .B (n_563), .CO (n_611), .S (n_564));
  OR2X1 g38932__7410(.A (n_1683), .B (n_1616), .Y (n_562));
  MX2X1 g38940__6417(.A (g336), .B (g1068), .S0 (n_1251), .Y (n_561));
  NOR2X1 g38916__5477(.A (g471), .B (n_509), .Y (n_560));
  MX2X1 g38959__2398(.A (g357), .B (g1089), .S0 (n_1251), .Y (n_559));
  OAI221X1 g38912__5107(.A0 (g1255), .A1 (n_481), .B0 (g1007), .B1
       (n_763), .C0 (n_480), .Y (n_558));
  OR2X1 g38911__6260(.A (n_464), .B (n_566), .Y (n_557));
  OR4X1 g38692__4319(.A (g396), .B (g426), .C (g401), .D (n_452), .Y
       (n_556));
  OR4X1 g38694__8428(.A (g496), .B (g486), .C (g501), .D (n_451), .Y
       (n_555));
  OR4X1 g38744__5526(.A (g1240), .B (g1292), .C (g1265), .D (n_442), .Y
       (n_554));
  CLKXOR2X1 g38748__6783(.A (g1864), .B (n_477), .Y (n_553));
  CLKXOR2X1 g38882__3680(.A (n_456), .B (n_431), .Y (n_552));
  CLKXOR2X1 g38876__1617(.A (g1419), .B (n_453), .Y (n_551));
  NOR3X1 g38871__2802(.A (g1415), .B (g1407), .C (n_444), .Y (n_550));
  SDFFX1 DFF_169_Q_reg(.CK (CK), .D (n_414), .SI (n_255), .SE (SE), .Q
       (g1411), .QN (n_27));
  NOR2X1 g38830__1705(.A (g1864), .B (n_478), .Y (n_615));
  INVX1 g38806(.A (n_549), .Y (n_612));
  AND3X2 g38878__5122(.A (n_1045), .B (n_548), .C (n_547), .Y (n_614));
  CLKAND2X2 g38917__8246(.A (g1900), .B (n_546), .Y (n_613));
  NAND2X1 g38920__7098(.A (n_545), .B (n_566), .Y (n_652));
  OR3X1 g38879__6131(.A (n_548), .B (n_1045), .C (n_544), .Y (n_648));
  NOR4X1 g38885__1881(.A (g1834), .B (g1840), .C (n_600), .D (n_523),
       .Y (n_734));
  SDFFX1 DFF_66_Q_reg(.CK (CK), .D (n_410), .SI (g327), .SE (SE), .Q
       (g1389), .QN (n_26));
  NOR4X1 g38887__5115(.A (g611), .B (g617), .C (n_467), .D (n_524), .Y
       (n_804));
  NAND2X1 g38888__7482(.A (g4175), .B (n_543), .Y (n_624));
  NAND2X1 g38925__4733(.A (g382), .B (n_462), .Y (n_1651));
  NAND2X1 g38926__6161(.A (g1231), .B (n_463), .Y (n_1360));
  SDFFX1 DFF_24_Q_reg(.CK (CK), .D (n_415), .SI (n_235), .SE (SE), .Q
       (g1424), .QN (n_25));
  SDFFX1 DFF_424_Q_reg(.CK (CK), .D (n_411), .SI (n_239), .SE (SE), .Q
       (g197), .QN (dft_sdo_23));
  INVX1 g38973(.A (n_541), .Y (n_542));
  MX2X1 g38941__9315(.A (g354), .B (g1086), .S0 (n_1251), .Y (n_540));
  MX2X1 g38944__9945(.A (g348), .B (g1080), .S0 (n_1251), .Y (n_539));
  NAND3X1 g38951__2883(.A (g471), .B (g466), .C (n_537), .Y (n_538));
  MX2X1 g38957__2346(.A (g345), .B (g1077), .S0 (n_1251), .Y (n_536));
  MX2X1 g38958__1666(.A (g366), .B (g1098), .S0 (n_1251), .Y (n_535));
  MX2X1 g38960__7410(.A (g339), .B (g1071), .S0 (n_1251), .Y (n_534));
  MX2X1 g38961__6417(.A (g363), .B (g1095), .S0 (n_1251), .Y (n_533));
  MX2X1 g38962__5477(.A (g351), .B (g1083), .S0 (n_1251), .Y (n_532));
  MX2X1 g38963__2398(.A (g342), .B (g1074), .S0 (n_1251), .Y (n_531));
  NAND2X1 g38987__5107(.A (n_1222), .B (g37), .Y (n_530));
  INVX1 g38975(.A (n_874), .Y (n_529));
  CLKINVX1 g38974(.A (n_859), .Y (n_528));
  MX2X1 g38939__6260(.A (g360), .B (g1092), .S0 (n_1251), .Y (n_527));
  AOI21X1 g38966__4319(.A0 (g1822), .A1 (n_429), .B0 (n_735), .Y
       (n_700));
  NOR2X1 g39073__8428(.A (g590), .B (n_1683), .Y (n_565));
  NOR3X1 g38969__5526(.A (g42), .B (n_526), .C (n_525), .Y (n_581));
  SDFFX1 DFF_220_Q_reg(.CK (CK), .D (n_423), .SI (n_77), .SE (SE), .Q
       (g166), .QN (n_23));
  SDFFX1 DFF_307_Q_reg(.CK (CK), .D (n_421), .SI (g1462), .SE (SE), .Q
       (g178), .QN (n_22));
  SDFFX1 DFF_97_Q_reg(.CK (CK), .D (n_416), .SI (n_249), .SE (SE), .Q
       (UNCONNECTED45), .QN (g1504));
  NAND2X1 g39007__6783(.A (g1718), .B (n_786), .Y (n_1119));
  SDFFX1 DFF_315_Q_reg(.CK (CK), .D (n_418), .SI (n_256), .SE (SE), .Q
       (g1520), .QN (n_21));
  SDFFX1 DFF_284_Q_reg(.CK (CK), .D (n_422), .SI (n_325), .SE (SE), .Q
       (UNCONNECTED46), .QN (g192));
  SDFFX1 DFF_118_Q_reg(.CK (CK), .D (n_413), .SI (g632), .SE (SE), .Q
       (g1415), .QN (n_20));
  NOR3X1 g38971__3680(.A (g591), .B (g611), .C (n_524), .Y (n_1113));
  SDFFX1 DFF_494_Q_reg(.CK (CK), .D (n_419), .SI (n_144), .SE (SE), .Q
       (g1515), .QN (dft_sdo_27));
  NOR3X1 g38970__1617(.A (g1814), .B (g1834), .C (n_523), .Y (n_1414));
  CLKINVX2 g38977(.A (n_1384), .Y (n_730));
  OR2X2 g39020__2802(.A (g30), .B (n_1222), .Y (n_1394));
  NOR2X1 g38902__1705(.A (n_399), .B (n_1686), .Y (n_522));
  NOR2X1 g38903__5122(.A (n_404), .B (n_1443), .Y (n_521));
  AOI21X1 g38905__8246(.A0 (n_408), .A1 (n_466), .B0 (n_1683), .Y
       (n_520));
  AOI21X1 g38906__7098(.A0 (n_518), .A1 (n_517), .B0 (g1690), .Y
       (n_519));
  AND2X1 g38910__6131(.A (n_443), .B (g1700), .Y (n_516));
  AOI21X1 g38942__1881(.A0 (g1250), .A1 (g1011), .B0 (n_441), .Y
       (n_515));
  NOR3X1 g38965__5115(.A (g471), .B (g466), .C (n_513), .Y (n_514));
  NAND3X1 g38967__7482(.A (g471), .B (n_511), .C (n_474), .Y (n_512));
  CLKINVX1 g38972(.A (n_509), .Y (n_510));
  INVX1 g38976(.A (n_566), .Y (n_508));
  NAND2X1 g38978__4733(.A (n_603), .B (n_524), .Y (n_507));
  AND2X1 g38979__6161(.A (n_523), .B (n_505), .Y (n_506));
  NAND2X1 g38981__9315(.A (g1657), .B (n_1251), .Y (n_504));
  NAND2X1 g38983__9945(.A (g1660), .B (n_1251), .Y (n_503));
  AND2X1 g38985__2883(.A (n_523), .B (g1857), .Y (n_502));
  NAND2X1 g38986__2346(.A (g639), .B (n_524), .Y (n_501));
  NOR2X1 g38990__1666(.A (n_459), .B (g32), .Y (n_500));
  NOR2X1 g38988__7410(.A (g456), .B (n_494), .Y (n_585));
  OR2X1 g38993__6417(.A (g611), .B (n_499), .Y (n_602));
  AND2X1 g38992__5477(.A (n_704), .B (n_472), .Y (n_579));
  NOR2X1 g38829__2398(.A (g646), .B (n_498), .Y (n_549));
  INVX1 g39026(.A (n_735), .Y (n_497));
  SDFFX1 DFF_275_Q_reg(.CK (CK), .D (n_436), .SI (n_257), .SE (SE), .Q
       (UNCONNECTED47), .QN (g1959));
  CLKINVX1 g39074(.A (g845), .Y (n_496));
  OR2X1 g39061__5107(.A (n_494), .B (n_487), .Y (n_495));
  OR2X1 g39046__6260(.A (n_513), .B (n_494), .Y (n_493));
  OAI21X1 g39044__4319(.A0 (g750), .A1 (n_427), .B0 (n_458), .Y
       (n_492));
  OAI21X1 g39043__8428(.A0 (g627), .A1 (n_426), .B0 (n_498), .Y
       (n_491));
  AOI21X1 g39031__5526(.A0 (g1781), .A1 (g1776), .B0 (n_430), .Y
       (n_490));
  CLKINVX1 g39025(.A (n_1117), .Y (n_489));
  INVX1 g39022(.A (n_488), .Y (n_1042));
  NOR2X1 g38994__6783(.A (g466), .B (n_487), .Y (n_541));
  NOR2X1 g38995__3680(.A (g1834), .B (n_486), .Y (n_601));
  NOR2X1 g38996__1617(.A (g1828), .B (n_701), .Y (n_583));
  NAND2X1 g39068__2802(.A (n_461), .B (n_485), .Y (n_873));
  NOR2X1 g39005__1705(.A (n_876), .B (n_525), .Y (n_874));
  NAND2X1 g39006__5122(.A (g1718), .B (n_1631), .Y (n_1259));
  NAND2X1 g39004__8246(.A (n_797), .B (n_485), .Y (n_859));
  NOR2X1 g39012__7098(.A (g1713), .B (n_626), .Y (n_686));
  INVX1 g39027(.A (n_971), .Y (n_968));
  NAND2X1 g39019__6131(.A (n_484), .B (n_1631), .Y (n_1586));
  NAND2X1 g39072__1881(.A (n_820), .B (n_626), .Y (n_900));
  NAND2X1 g39021__5115(.A (n_820), .B (n_1631), .Y (n_1384));
  ADDHX1 g38899__7482(.A (g4173), .B (g4174), .CO (n_543), .S (n_483));
  SDFFX1 DFF_445_Q_reg(.CK (CK), .D (g1854), .SI (n_229), .SE (SE), .Q
       (g7), .QN (n_18));
  CLKXOR2X1 g39059__4733(.A (g1011), .B (n_481), .Y (n_482));
  CLKXOR2X1 g39033__6161(.A (g1023), .B (n_752), .Y (n_480));
  NAND2X1 g38980(.A (g1727), .B (n_1379), .Y (n_479));
  INVX1 g38893(.A (n_477), .Y (n_478));
  AOI21X1 g38870(.A0 (g806), .A1 (g802), .B0 (n_563), .Y (n_476));
  NAND2X1 g38982(.A (g1724), .B (n_1379), .Y (n_475));
  SDFFX1 DFF_377_Q_reg(.CK (CK), .D (g101), .SI (n_36), .SE (SE), .Q
       (g2601), .QN (n_17));
  SDFFX1 DFF_100_Q_reg(.CK (CK), .D (g29), .SI (n_168), .SE (SE), .Q
       (g2604), .QN (n_16));
  MX2X1 g39049(.A (g546), .B (g1654), .S0 (n_1399), .Y (g6920));
  SDFFX1 DFF_62_Q_reg(.CK (CK), .D (g104), .SI (n_99), .SE (SE), .Q
       (g2602), .QN (n_15));
  NAND2X1 g38991(.A (g461), .B (n_474), .Y (n_509));
  SDFFX1 DFF_54_Q_reg(.CK (CK), .D (g1713), .SI (n_35), .SE (SE), .Q
       (g590), .QN (n_14));
  MX2X1 g39050(.A (g554), .B (g1657), .S0 (n_1399), .Y (g6926));
  SDFFX1 DFF_154_Q_reg(.CK (CK), .D (g103), .SI (g1397), .SE (SE), .Q
       (g2606), .QN (n_13));
  SDFFX1 DFF_343_Q_reg(.CK (CK), .D (g814), .SI (n_271), .SE (SE), .Q
       (g849), .QN (n_12));
  MX2X1 g39067(.A (g1811), .B (n_473), .S0 (g18), .Y (n_590));
  NOR3X1 g39063(.A (g591), .B (g599), .C (n_472), .Y (n_488));
  OAI22X1 g39047(.A0 (n_471), .A1 (g1690), .B0 (n_1411), .B1 (n_1399),
       .Y (g6949));
  NAND3X1 g39052(.A (n_470), .B (n_938), .C (n_469), .Y (n_582));
  NAND3X1 g39069(.A (g1828), .B (n_600), .C (n_468), .Y (n_1117));
  NOR3X1 g39071(.A (g617), .B (n_467), .C (n_629), .Y (n_971));
  NOR2X1 g39011(.A (g9), .B (n_466), .Y (n_1616));
  NOR2X1 g39018(.A (n_465), .B (n_464), .Y (n_566));
  SDFFX1 DFF_267_Q_reg(.CK (CK), .D (g636), .SI (n_367), .SE (SE), .Q
       (g8), .QN (n_11));
  CLKINVX1 g39024(.A (n_690), .Y (n_463));
  SDFFX1 DFF_295_Q_reg(.CK (CK), .D (g83), .SI (n_372), .SE (SE), .Q
       (g755), .QN (n_10));
  CLKINVX1 g39023(.A (n_1526), .Y (n_462));
  SDFFX1 DFF_55_Q_reg(.CK (CK), .D (g794), .SI (n_14), .SE (SE), .Q
       (g829), .QN (n_9));
  SDFFX1 DFF_248_Q_reg(.CK (CK), .D (g826), .SI (n_130), .SE (SE), .Q
       (g861), .QN (n_8));
  SDFFX1 DFF_412_Q_reg(.CK (CK), .D (g806), .SI (n_340), .SE (SE), .Q
       (g841), .QN (n_7));
  SDFFX1 DFF_338_Q_reg(.CK (CK), .D (g798), .SI (n_365), .SE (SE), .Q
       (g833), .QN (dft_sdo_18));
  SDFFX1 DFF_405_Q_reg(.CK (CK), .D (g818), .SI (dft_sdi_23), .SE (SE),
       .Q (g853), .QN (n_5));
  INVX1 g39075(.A (n_461), .Y (n_567));
  SDFFX1 DFF_309_Q_reg(.CK (CK), .D (g802), .SI (dft_sdi_17), .SE (SE),
       .Q (g837), .QN (n_4));
  SDFFX1 DFF_150_Q_reg(.CK (CK), .D (g28), .SI (n_82), .SE (SE), .Q
       (g2603), .QN (n_3));
  MX2X1 g39051(.A (g557), .B (g1660), .S0 (n_1399), .Y (g6932));
  SDFFX1 DFF_367_Q_reg(.CK (CK), .D (g822), .SI (n_381), .SE (SE), .Q
       (g857), .QN (n_2));
  SDFFX1 DFF_433_Q_reg(.CK (CK), .D (g810), .SI (n_270), .SE (SE), .Q
       (g845), .QN (n_1));
  NOR3X1 g39056(.A (n_469), .B (n_470), .C (n_938), .Y (n_546));
  MX2X1 g39048(.A (g560), .B (g1663), .S0 (n_1399), .Y (g6942));
  SDFFX1 DFF_129_Q_reg(.CK (CK), .D (g102), .SI (dft_sdi_7), .SE (SE),
       .Q (g2605), .QN (n_0));
  CLKINVX2 g39076(.A (n_626), .Y (n_631));
  NOR3X1 g39070(.A (g1840), .B (n_600), .C (n_460), .Y (n_735));
  CLKINVX2 g39079(.A (n_1251), .Y (n_786));
  INVX1 g39077(.A (n_459), .Y (n_1222));
  CLKINVX2 g39078(.A (n_458), .Y (n_1669));
  CLKINVX2 g39119(.A (n_1631), .Y (n_1149));
  CLKXOR2X1 g39038(.A (g521), .B (g525), .Y (n_457));
  CLKXOR2X1 g39058(.A (g1003), .B (g999), .Y (n_456));
  CLKXOR2X1 g39035(.A (g1235), .B (g991), .Y (n_455));
  AND3X2 g39036(.A (g744), .B (g743), .C (g109), .Y (g5659));
  CLKXOR2X1 g39053(.A (g1415), .B (g1515), .Y (n_453));
  OR4X1 g38901(.A (g448), .B (g452), .C (g440), .D (g444), .Y (n_452));
  OR4X1 g38904(.A (g530), .B (g538), .C (g534), .D (g542), .Y (n_451));
  CLKXOR2X1 g39045(.A (g1015), .B (g1019), .Y (n_450));
  CLKXOR2X1 g39029(.A (g1845), .B (g1861), .Y (n_449));
  CLKXOR2X1 g39030(.A (g1260), .B (g1019), .Y (n_448));
  CLKXOR2X1 g39032(.A (g1265), .B (g1015), .Y (n_447));
  CLKXOR2X1 g39037(.A (g1240), .B (g1003), .Y (n_446));
  AND3X2 g39034(.A (g742), .B (g741), .C (g109), .Y (g5658));
  NAND3X1 g39039(.A (g1436), .B (g1424), .C (g1444), .Y (n_444));
  CLKXOR2X1 g39040(.A (g1707), .B (g1690), .Y (n_443));
  OR3X1 g39041(.A (g1300), .B (g1304), .C (g1296), .Y (n_442));
  CLKXOR2X1 g39042(.A (g1245), .B (g999), .Y (n_441));
  NOR2X1 g39140(.A (n_1359), .B (n_1399), .Y (g6955));
  NAND3X1 g39057(.A (g658), .B (g668), .C (g677), .Y (n_544));
  NOR3X1 g39054(.A (g658), .B (g668), .C (g677), .Y (n_547));
  NAND3X1 g39055(.A (g45), .B (g44), .C (g43), .Y (n_887));
  CLKINVX1 g39118(.A (n_513), .Y (n_537));
  NAND2X1 g39107(.A (g44), .B (n_428), .Y (n_525));
  NAND2X1 g39104(.A (g466), .B (n_393), .Y (n_494));
  NOR2X1 g39111(.A (n_425), .B (g1703), .Y (n_626));
  OR2X1 g39085(.A (g1771), .B (n_439), .Y (n_440));
  INVX1 g39117(.A (n_1675), .Y (n_438));
  NOR2X1 g39084(.A (n_436), .B (g1707), .Y (n_437));
  INVX1 g39115(.A (n_434), .Y (n_435));
  NOR2X1 g39128(.A (n_1683), .B (n_432), .Y (n_433));
  CLKXOR2X1 g39060(.A (g995), .B (g991), .Y (n_431));
  CLKINVX1 g39116(.A (n_464), .Y (n_430));
  NAND2X1 g39100(.A (g456), .B (n_511), .Y (n_487));
  NOR2X1 g39112(.A (g31), .B (n_829), .Y (n_459));
  NOR2X1 g39137(.A (n_467), .B (n_472), .Y (n_499));
  NOR2X1 g39143(.A (n_600), .B (n_429), .Y (n_486));
  NOR2X1 g39108(.A (g44), .B (n_428), .Y (n_461));
  NOR2X1 g39102(.A (g1861), .B (n_407), .Y (n_477));
  NAND2X1 g39113(.A (g750), .B (n_427), .Y (n_458));
  NOR2X1 g39105(.A (g43), .B (n_888), .Y (n_485));
  NAND2X1 g39106(.A (g627), .B (n_426), .Y (n_498));
  NAND3X1 g39062(.A (g971), .B (g976), .C (g981), .Y (n_1686));
  NAND3X1 g39064(.A (g1336), .B (g1346), .C (g1341), .Y (n_1443));
  NAND3X1 g39065(.A (g378), .B (g369), .C (g374), .Y (n_1526));
  NAND3X1 g39066(.A (g1227), .B (g1218), .C (g1223), .Y (n_690));
  NOR2X1 g39109(.A (g591), .B (n_580), .Y (n_704));
  NAND2X1 g39149(.A (n_580), .B (n_472), .Y (n_524));
  NAND2X1 g39110(.A (g1822), .B (n_600), .Y (n_701));
  NAND2X1 g39150(.A (n_429), .B (n_468), .Y (n_523));
  NAND2X1 g39114(.A (n_425), .B (g1703), .Y (n_1251));
  CLKAND2X2 g39154(.A (n_425), .B (n_391), .Y (n_1631));
  NAND2X1 g39123(.A (g822), .B (g818), .Y (n_424));
  AND2X1 g39122(.A (g143), .B (g109), .Y (n_423));
  AND2X1 g39129(.A (g1389), .B (g109), .Y (n_422));
  AND2X1 g39124(.A (g148), .B (g109), .Y (n_421));
  NOR2X1 g39125(.A (g1766), .B (g1713), .Y (n_420));
  AND2X1 g39135(.A (g1419), .B (g109), .Y (n_419));
  AND2X1 g39120(.A (g1515), .B (g109), .Y (n_418));
  NOR2X1 g39130(.A (g794), .B (g798), .Y (n_417));
  AND2X1 g39121(.A (g1499), .B (g109), .Y (n_416));
  AND2X1 g39133(.A (g1407), .B (g109), .Y (n_415));
  AND2X1 g39126(.A (g1424), .B (g109), .Y (n_414));
  NOR2X1 g39139(.A (g466), .B (g456), .Y (n_474));
  NAND2X1 g39144(.A (g814), .B (g810), .Y (n_594));
  NAND2X1 g39141(.A (g1786), .B (g1791), .Y (n_518));
  AND2X1 g39131(.A (g1520), .B (g109), .Y (n_413));
  OR2X1 g39134(.A (g48), .B (g30), .Y (n_412));
  AND2X1 g39132(.A (g1374), .B (g109), .Y (n_411));
  AND2X1 g39127(.A (g197), .B (g109), .Y (n_410));
  NAND2X1 g39142(.A (g109), .B (g1453), .Y (n_434));
  NAND2X1 g39138(.A (g18), .B (g115), .Y (n_466));
  NAND2X1 g39136(.A (g1801), .B (g1796), .Y (n_517));
  NOR2X1 g39147(.A (g45), .B (g44), .Y (n_797));
  NAND2X1 g39148(.A (g109), .B (g201), .Y (n_1675));
  CLKAND2X2 g39151(.A (g794), .B (g798), .Y (n_563));
  NAND2X1 g39145(.A (g1766), .B (g1771), .Y (n_464));
  NAND2X1 g39146(.A (g43), .B (g42), .Y (n_876));
  NAND2X1 g39152(.A (g456), .B (g461), .Y (n_513));
  NAND2X1 g39153(.A (g1696), .B (g1703), .Y (n_1379));
  CLKINVX1 g39219(.A (g554), .Y (n_409));
  CLKINVX1 g39161(.A (g9), .Y (n_408));
  INVX1 g39166(.A (g1845), .Y (n_407));
  CLKINVX1 g39206(.A (g881), .Y (n_406));
  CLKINVX1 g39171(.A (g677), .Y (n_405));
  CLKINVX1 g39226(.A (g1351), .Y (n_404));
  INVX1 g39207(.A (g23), .Y (g3327));
  INVX1 g39176(.A (g4176), .Y (n_402));
  CLKINVX1 g39173(.A (g374), .Y (n_401));
  INVX1 g39177(.A (g826), .Y (n_400));
  CLKINVX1 g39222(.A (g986), .Y (n_399));
  CLKINVX1 g39163(.A (g1304), .Y (n_398));
  CLKINVX1 g39210(.A (g1621), .Y (n_397));
  CLKINVX1 g39181(.A (g1245), .Y (n_754));
  INVX1 g39191(.A (g1766), .Y (n_439));
  CLKINVX2 g39156(.A (g1666), .Y (n_471));
  CLKINVX1 g39184(.A (g426), .Y (n_1661));
  INVX1 g39239(.A (g1900), .Y (n_932));
  CLKINVX2 g39217(.A (g4172), .Y (n_427));
  CLKINVX2 g39162(.A (g546), .Y (n_1624));
  INVX1 g39215(.A (g201), .Y (n_473));
  CLKINVX1 g39174(.A (g1700), .Y (n_436));
  INVX1 g39195(.A (g668), .Y (n_1043));
  CLKINVX1 g39180(.A (g1235), .Y (n_757));
  CLKINVX2 g39159(.A (g575), .Y (n_1083));
  CLKINVX1 g39230(.A (g1265), .Y (n_779));
  CLKINVX1 g39231(.A (g1240), .Y (n_758));
  CLKINVX2 g39167(.A (g1411), .Y (n_432));
  INVX1 g39242(.A (g1834), .Y (n_460));
  CLKINVX1 g39198(.A (g45), .Y (n_428));
  INVX1 g39183(.A (g1801), .Y (n_788));
  INVX1 g39213(.A (g4), .Y (n_1291));
  CLKINVX2 g39218(.A (g563), .Y (n_1411));
  CLKINVX2 g39193(.A (g1872), .Y (n_470));
  INVX2 g39244(.A (g1822), .Y (n_468));
  CLKINVX1 g39188(.A (g658), .Y (n_904));
  CLKINVX2 g39238(.A (g1270), .Y (n_752));
  CLKINVX2 g39202(.A (g591), .Y (n_467));
  CLKINVX2 g39241(.A (g611), .Y (n_629));
  CLKINVX2 g39197(.A (g722), .Y (n_1046));
  CLKINVX2 g39240(.A (g1918), .Y (n_935));
  INVX1 g39170(.A (g713), .Y (n_688));
  INVX2 g39200(.A (g605), .Y (n_472));
  CLKINVX2 g39201(.A (g1814), .Y (n_600));
  CLKINVX2 g39247(.A (g1713), .Y (n_820));
  CLKINVX2 g39248(.A (g1690), .Y (n_1399));
  INVX2 g39249(.A (g18), .Y (n_1595));
  INVX2 g39250(.A (g109), .Y (n_1683));
  INVX1 g39179(.A (g511), .Y (n_396));
  INVX1 g39155(.A (g950), .Y (n_395));
  INVX1 g39209(.A (g1394), .Y (n_394));
  CLKINVX2 g39246(.A (g471), .Y (n_393));
  CLKINVX1 g39224(.A (g1796), .Y (n_392));
  CLKINVX2 g39223(.A (g1703), .Y (n_391));
  INVX1 g39229(.A (g4178), .Y (n_390));
  CLKINVX1 g39212(.A (g1092), .Y (n_389));
  CLKINVX1 g39160(.A (g105), .Y (n_388));
  CLKINVX1 g39175(.A (g1403), .Y (n_387));
  CLKINVX1 g39228(.A (g1223), .Y (n_386));
  CLKINVX1 g39169(.A (g1786), .Y (n_385));
  CLKINVX1 g39233(.A (g1260), .Y (n_765));
  INVX1 g39220(.A (g560), .Y (n_1478));
  CLKINVX2 g39157(.A (g1868), .Y (n_616));
  CLKINVX1 g39234(.A (g1857), .Y (n_505));
  INVX1 g39168(.A (g1776), .Y (n_465));
  CLKINVX2 g39211(.A (g654), .Y (n_683));
  CLKINVX1 g39196(.A (g1781), .Y (n_545));
  CLKINVX1 g39186(.A (g1718), .Y (n_484));
  INVX1 g39164(.A (g4181), .Y (n_951));
  CLKINVX2 g39208(.A (g643), .Y (n_426));
  INVX1 g39194(.A (g1791), .Y (n_692));
  CLKINVX1 g39214(.A (g572), .Y (n_1244));
  CLKINVX2 g39158(.A (g569), .Y (n_1299));
  CLKINVX2 g39182(.A (g481), .Y (n_650));
  CLKINVX1 g39203(.A (g43), .Y (n_526));
  INVX1 g39221(.A (g1945), .Y (n_800));
  INVX1 g39227(.A (g1927), .Y (n_717));
  CLKINVX2 g39185(.A (g1007), .Y (n_481));
  CLKINVX1 g39187(.A (g1250), .Y (n_755));
  CLKINVX1 g39216(.A (g557), .Y (n_1563));
  CLKINVX2 g39165(.A (g566), .Y (n_1359));
  INVX1 g39172(.A (g731), .Y (n_776));
  INVX2 g39199(.A (g1828), .Y (n_429));
  CLKINVX1 g39205(.A (g48), .Y (n_829));
  INVX1 g39235(.A (g704), .Y (n_649));
  CLKINVX2 g39243(.A (g461), .Y (n_511));
  CLKINVX2 g39236(.A (g1255), .Y (n_763));
  CLKINVX2 g39190(.A (g1936), .Y (n_937));
  CLKINVX1 g39232(.A (g1696), .Y (n_425));
  INVX1 g39225(.A (g695), .Y (n_548));
  CLKINVX2 g39178(.A (g1891), .Y (n_469));
  CLKINVX1 g39204(.A (g42), .Y (n_888));
  CLKINVX2 g39237(.A (g639), .Y (n_603));
  INVX2 g39192(.A (g1882), .Y (n_938));
  CLKINVX2 g39189(.A (g686), .Y (n_1045));
  CLKINVX2 g39245(.A (g599), .Y (n_580));
  XNOR2X1 g2(.A (g976), .B (n_1687), .Y (n_1731));
  INVX1 g3(.A (n_1732), .Y (n_1733));
  MX2X1 g39685(.A (n_1658), .B (n_1655), .S0 (n_1338), .Y (n_1732));
  XNOR2X1 g39686(.A (g153), .B (n_1628), .Y (n_1734));
  CLKXOR2X1 g39687(.A (g162), .B (n_1573), .Y (n_1735));
  CLKXOR2X1 g39688(.A (g174), .B (n_1482), .Y (n_1736));
  XNOR2X1 g39689(.A (g1341), .B (n_1455), .Y (n_1737));
  XNOR2X1 g39690(.A (g170), .B (n_1416), .Y (n_1738));
  CLKXOR2X1 g39691(.A (g127), .B (n_1366), .Y (n_1739));
  XNOR2X1 g39692(.A (g131), .B (n_1306), .Y (n_1740));
  CLKXOR2X1 g39693(.A (g135), .B (n_1247), .Y (n_1741));
  XNOR2X1 g39694(.A (g139), .B (n_1111), .Y (n_1742));
endmodule

